`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FKyl7WebfaCvtrIdsiNIsKAJHMSc1b85D7Dqp+mvmI2Oy5AxMtjaa10KVNe2hsR1phi85jax4+/+
i5Ie2C5e+w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Etda3DA4SBU8KpHadhe1aXzCa2697lfsClupRip/dJk4Op6J7K6PJTHrHSCU7Tj7RX0EFcP4bzQW
xQTG6xveUqXfaPBigSeIO2vG8z75o6PDp/wIE/rT0W4KsB3v6DxLiJyibYl6Vcu15jK9VeCHtRmB
bLBgWsFP/E1/47P4vRg=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Du3bkjkphrTJhJxNd71iXfb4lQ087sdSdm98c0YeW5PUqriRhHjYv6e3LN4EcDSqM68XOiMTYUJI
gpomXpPyCpPibqrDZZsLTutaLGd0hQSKrfCXg2sL7aAhZyiKFQCt4+lWenWr2wM/+XAo2AZD2yWA
vDffpMh6OOWo72zEQdQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VkwBgHuAYuNsjW85cJFAwFYSe3fb1ScFnAGcE0Ek/zbD1F+WMDmKWXaCwrts7qx9LTBsAUWqFSOz
WYprRa1T5j6uPOc4JLyrDFLTVaAnGHsAXJpusv49XfG6eWrjPI8+fQsWRKGRJ8tvsdndbbDHbFRu
PlR5HQWuXAfqkXb+dp6zzdOQdUahOaQr7nFpYsTr4FxkbVQvmCt8grUhAJmHhK4nyLE+g1noXq3Q
mlNWvntZwf6h0AON1yxD9GyLMkUg+EWZ/U92yuo21KE7dwVdgPovYyDZd4NStgVJ+ixmAjK+xhfK
VH9hHKzeHaiLkym6g7HLpJZ/TzBvG6bt2gRfMQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VLTWuI7riGPMgTH6sPnohEwGDWG9kiM/HIkMiWt1wAHbn68V+36cwvFcqhH51ur6fors0ZplVg/p
rhqRdrdjmEDsq7/wDF1tfnnp5r5SF4TSRNO6HnasRKbYaMjHB70qWLKvZSVUPYYNmVUIodMAorta
5meyAj0qbVPkiCJ5UUg9AXBXDj+IcU2VbV1oMrRVzI4HaIrpTbgVPaViNXh3pLCQHLEB1FbnkFJ3
5CUWSufH7e8RfKd658XHnntcUuAX20B0gvJ875n3qVMr2irr/zISF75DeOdvYVrn0ZqUZgpWSvGB
bSlvgKC/dV+kuOw2raFhY1VCmcSkPZ5dprN9/g==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HDrBYpliRrBIBPVo8k/EgNJjvaTocIUlpspjLQIJDo3w+nSeWzXL01GIojcxHLBypyhQ1YXOYQTO
PJN6T9UkDvu/4L87I5lnu7f1pTGuE/ri9irkozP6M4Odtsxws7hnWde78sA5V4gV8u2nmPGlRX+s
PlnMABrZ2EKLMNXWYwtFQpMXGCgyfW26y5lhMce/IKJaee4hbeD5PDJbGfbQbyhIU9TpZthaGQsZ
UcROvfYe6wJUAnoRw9qtReAXYWAKDoktAsVPYL43ump3nBdNvJKVcLJd2gD8q9HWHBWDLaUAhba3
nRh8Pi8N3TxwfwBFloS3kWk+PxYhRkvJvQBIoQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 211040)
`protect data_block
o4tITWbOoysjjWjH/Uupk6FqrG7Q50YWdXqT0gkhDNkRTgaB0v1ol6bOsQiELK2Nxg32iZRiDlBI
ZXGt+9GlsO1T0Cc/nkxnq/PPoWk/264tTimHc2x3lrGmkDXjd2ZH9dx+yXmsMyq9MbQWqCIWOm/E
rgASaINGiTBT7JE0+N+DB3RCCWEIaed2P+7yf4vFpo/vEzNpA7z74qRrHJT3WwOgIPJV8755kDfM
NV5nfKWL30bAGEk1l0wki5hfas7ye6op5+iLOH7BVr/awuJCQqmagvFqZuOmYgFMR5PLclVdg+O8
SRoahgTkwFTWQIE0VFprPsphgtBjDkmfQNWlbbPhvLKYDf7a8HBhzHuOCYHnPkhNVZBMAsWg4ueN
7/z54Pt+4lQuG3bIoq77mT4uu3uskQdpiYFzSumfVfr5M0+R6aaEpeM1MVQ9EI+jduWw1okV3QnE
d9mHYuMJMixgDMx3ruhf4mYrfF3dCaGqbJr0meefS6kWWwCg980yt3ZxA8OuIrkxNWfHar8TTn/A
uYN3iC+kumzni8GD26S8GASlpnirJ5LPEJgqUx4L6jiAClOmst4/nkZD2YMtD/W7spaSbZ+jJg9b
7/jsIYkC6nnPt4cvzY6q9SRv2q2Fm9ppOuX4P0m7nS9NJUCghzoKH6WTThWdoN/vjXP4dusPF9zt
EdtLiPiGhLENSQdXqVjasBTmEpnNvxBmxMJL80N+oSAK5bR8dQA4sE/5lkVQBDJmkJ7xKETM5sKb
3hdm0v9lq7A2eMU5GvOpFLhBos5EV1rzsBtRglD3RNkWlgxNth4ZBrFM9adMBE9d6mYvGknBtN3K
2HxXiTxhnBkEvxA4nU7QHW8rpJ13YSNitUQouUhSvwMTaa7sROdnR60SlJIzUM5rFd1sEqq8w81I
jnH1p0GvIutk/9bDpeEZ9BGNsAov/jFdyOOCUb1scinL4e9lhEXyvuWrRYWvsG/HaesEVpDvAtoy
i0Bn/y7mR4A0tB6F5SOpSItshXiwpNCoKeN6Aw9xdDgFMvw4FyPyx9V+nyIowgAU0gmvLkMY9zT6
ubeypiUGBancxfSzx0TEWAFCPevj59HY0Ym5ChCu+aBllMpea1fC1yGUsdCwCVaunnwvpH06YYBQ
H9cvLpuYwVTgDIx4qMmp/whcCbbThFGlyaaj90Jh2OV58i7d29jdSS+zS3+bGzkHAI2jzBd+ARgR
VZiBUTFnOxCsSGmOxosUbIXy5YCl5DsFAxblltk3yRGP+BkCX7qpeEofPPxHzD9/7Da4UbUAxE+F
L9jpJBkqRT7c0aTkMUFNhzIFlrpEfTM+T34wdejwdBnR+icb8969YXQsx6HLI7okYuzrfBq4gD9e
ghxRFku9JaAQEBVAZe90XFMMgPS6YeTcxW9fNkc4JttyxJYrVfb2PCJExrnOZztZqRSglq272g8Y
ayrDStFTqwvR62ZzDyPwdo6jKtNboxoLA8FatzOe369SQZvduPwM+DO1o4ecOdHVF3OMM7RLXVIj
erU/FmZysaogOMzw58trWnxZLtLZuOJTm7Vm0GBOE/cpxf76bILp4TCB4XaB+0imA5J50mDvzFdu
bSnq83uku4a8rX7RU2HJBhWBve/AZnh5Axxob4QegdCN9qBeHspQw3BP6IJtBg3yQZL/c9GZv4Ts
LsY3yoRxTTxvehEhw/UoGnG4q2SxAgh5gFTn3WkAk1qTcSKpoN8EfGUMiT9aQC1QeBQ50kNCq+7K
ZeU+W8Afhpe2pHsFzGnLeG6Q1qsnklgf2WgPI/56Tq12BhQv6400DtZ14FeCYIC3u9P03yq1kQIl
Mlw/XPlz+2y6autS84lAe/1iyRo9Vx6Mez92TliKUvrCk41XFAmSJcWOI43hHfbosVWThsqrmwQQ
EYKJaiCrRUEJv88H+f6O0jdsc9T2q9UvSKKc+fkFnNx/2NTtHJivASj/45aS0K0EtxTpgwI7CSgX
poLbg8fbKmaU8hT34AaaiE7bmXJaF0+Nn5E3/sAfK8nfje1favYUwfrJRvhaXXrOdrAfPdEQ1R9n
mJq/iHP9NK35KfWs07jPJ0OzIynaSoAsF844C9ANeHOPtP2kzpI/YZNDC1Q9U6WeQirRrITGFikV
xcbLoXBSnBbms4ZjTUE6TQmIfv2n/ilLrO/9WFTazoHSJmpH8e9U5nFTYrpBIMeEcjlpjUJSgDk6
NKiHxD1Uv8AszK79lVQjJAHssmxu/X3DvmaFTONgwdYwDz9+dtTNHOMXQaOqKyUe7ue7zAQGdCII
5SLu01rdiu/LMXpLEYEnGuwHp4r1dbvLoPJWp0vDz971/yhOkyfgCqPPT6OVInXXKDlv+ioG+IPy
y+gnp2IMns3oDeaxBMyWbe7cV7FnVnQFpD+vSJtoj4ge7eJ+3v1vpCz6zQzNJlp4VvfliQByIXLA
fXzAG/m6LrabJm9iKMDSE4iJJ/iPyGrKnDP4kd9A+LEBkTFEjFKMJ8Qz3BB8sJAc0iB76n8lGl3h
+56voIKmN7P2aVO95NT9ZdFvD2dWLuB5UoyEfoaQDICPAwSDm9eT5YCkMIbV7WbFrM9BxdcckZyH
uX4JgSDpNgIaBWeUXiWnh6AT+RVZchBGFTTCcQtAOWR7QdGe+hOoXh8LFeNxKyfKfGhIFcGeeIsc
lfVR89Dk7JCUQuL2ywMzynbzwy1RLGX035L/m4aG+9vC7X9NmZe2PnPowSImhH4M0umdpPlPZiGm
9mi+aZ5oP6enbr27IUmIE/9M+OirR/6cvZ/0y33utE0aowe5Q3ZbSl25Ssl7n7PX1eS9cf4W7Njs
Qk8CDsRbek0iaMwe9Vb8UYFzeapXstNyKjCGq5E3VoOlpy5sSXApSOHS239ATVLE1PWF1LJrHRO+
LhC3Dd5kjHV1CvnAUMpXQuffUuSIt4p16Z1xiZmr2qe7jBWcVjxpuk2J0Dn7LhJ/Hkq0ykqYI5zI
tjkNGgAInB8kwZyvEHUpsuQS2sSJM1T7WxpfOi9aRUv0bKSirr+7ohufR7vHJFyAbleYA7J8D5ug
Vo7x+HCrV3roXnttDoh8RhxfhlUrLmw1hwbJUKYe7AfBnubJKEjXZuVkOcpj/2VU7eS3e9vFe8Mb
EtN39acLIWNXqCbjqBZWVxHvGU1Ezm7N4TP8c7s/Y31dWpYSoR8N6oofdzRGrXsGV9hbv6O04LDk
TgENuc4gHnU6aXSaq9fr0fG3qIWFYrQ3WpFrEGSI6zm0DWflm1H2KGr2p4FL6GydYjox9Yq56b3G
aK65E+p3Cr0mYa1RqLSnsn0VAIRhEQmXzCHvspMn1yTNN2WfKUVlF4Gk7toCYlvgCO68SiBt+g3z
u/yLS5e+5nbPr2Gb795fHxmR11Tz+1w6O/4Wh5mMUjJx7Su3KWoV9PLX/iwSQwqzdVyv18FUfkMm
yT2Xb6Xo3iTNVCHSG9ASkN2EpSa03yoP48e7MpozA6w5/cHyBzywHORdCN2QpKAGjpU2QOkS5Hc1
9VxHjZX2qQu+mw3+cGeU+SLI+mkkvqnfd5zVae2bSfnfHLzTxqgImfK+D76o3RAH5NgwOTXHykkL
+setSuAEWIHEqYJBf5hJ9+WXZH+O2PVUiMPr3bIZG+Ea9Rd/QCBHNYDl81q1PHgxeQb4gD5oqOQC
Ud/VvozP1us2Js3KYQdzYbaT9B+oNckQH3adHzxw/Nof3YVKKOyKA8wUkTpwTuiUqX07sxJjk3Xa
bth1G/TW6TcXjj5Aof6PQWOvKPrHEfnwoYp5YRuIE3Fg+1DgGShkm39qiwgz4IbSNnSjMNE5Ph/Y
Z/lhOz7Qi6qpV9/bs+seHScOO3J4K4ekxU2ioq/1TCSBFOCCSW2ilU70Uqdakhfzb2EffwsNFiY3
wa0wkWnPLsejuzXx7TnaY+t6h8lxolvzM73dZfaJK9HvP8TKM7NsJI73/bZjKV7DY5UDjczjmCry
PdZs+oj3dYXZzVej8TV9M/DZnmG713phIpU87cruf3p65EL5Re0CDotNud2ileBljE0PcGoFqcru
7Y95ipSIeHAjWsmJaCi4UTnfOUxy0QD+Ca0wFJ9fZLJ1oNLiRFOLoucs7rzxV/72aBzdsp2Ece3W
Gp5t6OBcjVbpYIlrDdbon6+Gt0hRYRzJ9hlROV1v9iM2K7hmInWsVN6ch8ExzYo+x1REXjwqHyAC
Nr9jJZXTZfbhZd1sL2RoHwU+4E4I1hBiC5VFmZKrmNwb2LTJKhbP3UNeSFcujgg089c5SuYdPsP2
FDI5XYi+lPs1c7/zhrgLoDnc31oB/HKmFIAIgxBE5eDb9l3NBz5xEv/bNbRWS/7xrJq0FBCMdqPs
w+2rodNi+0frO6yO4ZcH0Zx8DwKXlizt/TsGizvGylJvTEX4UMDhToxnQ4ATLXlaxRhf9eWTs9YC
7ESuQRRBIHwmQVc00dAD0z/R7HgVxxfI8TwxG+RFXgme20sE614Nne/7RgzzfYJVMFFBrEKemdbH
IwGWITtxqk5RHa/N2M6OKXuZ2Eo9Q42MwFeHyrUQ+2TF+g32LQN/z1nyiR8Ivu1px5UCNoISKwk1
lI2MiJPXISgBjRlZNqnqKsodI6SPJrHYHaeGl5knSuj5/uY7CzxMfWtAjV2llurqSQCp82mH8NvJ
LuXtwu0qoDvwCkivFMR9fGNSC8iJqYxnWtHI3bIpsPIxYFv6jJ5l/gB2E5tzNwI/DOUr1DHPLpBo
cUbJkKTnuI2GZ24pC3NKNGhQd3Q5BKn8zPiOFaaVRnA/ksr4bI+fvApMutSQx63DUTW2mD8Fw8/a
Q7aSLIlEx72+MvwjT48RkWT7FBJLg/zhCami7oGtHtcRYFIE+viHVak8Z6jhQ9y/Wh1hYrhmK070
/k2wSNuzaZTkTRS58qVxQgnFNOHR9aoT+IPO9ObgE3QSMsvoXPUq5aJzR2rwoXsG4yW8uKSirMlo
4xE+X50ICeIOoYVwo/d+rToWeoDJGHGSVCKB8nB0A+Rd1ay0m8a9oWIZ+26fc+6GW88n3hMx+5lz
PiXkubeGc8pTpiWBbaz5s+WoOduavFGp54Qu5cD2cYcqb2KA3N3yqLnk++9P5vpE+OPoSSx1xKTg
M3TBr62doEe041YWvaXx1/ryApKy8ic/juLH+YqnxMGeS8yIcCS5kf4EYFjkZcaoxswbBkaGlAPt
YombQrwYAPpU0s0mSgUtVLDNSbeYoORH5Ay2dQBZbZA34Pihn3EGXPaLse44rFCwbgIvJiQHBlqB
mhb589bQB7/Jszqn2Y0Dntzq0WI7rVnRSsN6WTCSKR230kumJwvxq7VyeUPt7t7WoUt9GL2VY25Q
A1xDCmEIL2MGafW/QMI7D3sJBLqCVd0A1j1Wju6KsGJjSwHyvGhln2iCI7sSLpv7F9ExSi3lD//Y
yu0yRKrjYFPrHLUq1pV/WZryt/CY/9mCzCEQrIA0DeafwMe+E3PBDGLFcn4aiAgfp9tfTTPzUGfN
Cn9+IWwKZKO49DOcloYJDeCXXjtzJjj8cTjSddw/3LnWUP1BXulZ6kjsya8Vxtqwk3JkDKMQBWhs
RNm6AF8T5pElrRogoN+3x8oFlb0lOkk8CKrTFeGWOTsKI3YtR9SQzmx7pHYKWfWdOCGXZa6QHSGM
WNEF4IxBmtOzRxMYvAHukQRYBygTndxlzBHPfpGwqxGrx6+8gkOVC9pG/BycTIpl10P7iCpdAltN
ZtuzrIF8vkheFOx4MK5ptdGbRFwW8OZwWBwwKGbqtDcOvuCgblL5nLanvEOXEvzWtLdJjeg7jbiO
dzIM2q13JHhlEpi+3KdnYkm38XwXO0wFpxjzf34vIAW++EPuWSPJOaAZAiyCduMe+KQ3uI6hNzYf
Lkpx27n6YNDn0686TmYoBudty9qj7JanXK/tqLL74TlHdNGbr1LnMjY5PoXP+H9cRm2GlSN9JOIB
BZMcDNurUmXmzNeNRVeiEBtEdYJoqYdRJD/8zPZDeGtRnNCxulQiTXGM36NLPs0/+2HzpKOe8ekp
1zCSDML1MYr+KYsDOVBTPmHiu9s4akxNf38hSIotjuVcBzJLlfSLlmOExV8D7hJThY25MhHONHZ1
6W2uy0jH7/HVt2a4JP5+IGxWivJEkLmsPciqY2gJk/5bRDvGLnYWu1Wkf+pvmjcxyQ4/C6mg1MzC
N06cdBm3INQzkCrylbBqQyosbFWLloZyrgWNoDfg2cPw+JIW7xAzyKFNoGX0qGgGQdXdLodK7jD4
2a26IXgByxzMbt4bGlrjgdVBOaVgeIWfMMl0G2ZdqJRw2W6vDseaPFuRxRJaXUi3WsP/QevHIMj0
kQ/iKjUTjtw5yR77w0KVXkpG5GOSx0hZg1yx65TCThlBDrmhU2GhJFVdAPPFu4PMDQKvYI3bPYio
/oaTd3EpP5IsK9uBa7pyh6HGIjNDvJdNo2SmlztQwm6+vNB/Npt9JTD9iahssE4pURMhcsSC4XBq
4MMiBPf4wjEAy3/mtlCHkAsxG78ETWyh3mgmkRuVk3Pxnc9981dqXb+QmyPR1KNxxseQzS6Rq3Ot
xa/yWbsEUVT1OvJj4wkt0acxASE/t80QkhsB0IQ5Lkp8mA9I961REZUX7UjYgricV1cM/UYaerml
6aN9L5NX9cbmqgUtpzFehED7etl+xDodN9vqXiCyz6zhAjHVp3wqaOsLkKcETEaJSjJbTuEH+Ki1
ew4oCJnNUGudxaE905lANKPRPkFGDEZWzyY5/bmi40rn6ukgOhAYDaulPrFbnz+kvbLn3y9dBS8z
hTmSKUCJ2kTFRYz7FUyOxJ2zKfVUvlNQvo+rZ5RF7BmexMabCE6prlzUkpvCxGlVjD6/XmPVuzq9
CnxI9Cdl1N4TJoAMNO8HjQPZj5I4Eqrpk/Ge02OjY6/HIYT7+yRNJkJa6vd5iWZz/Ng8AIXMUczO
U0LSFzkVgKcezr7aepare19yKdqZkIvg8qlzKd7uZ8ZH0iH93z2cA5REAUDHmDfxUPXZkbe0VzWW
IlTSegHk5XfsC3VKkt6DrgGH1/GEQ9gxBlrVyzshSUyddmw5mTeuBCEoIq5xYvVDHhjAvhkHVLNJ
wWZZoY1Vpdjv6E12JLEj/p++9GDt2OGI5MldKL4cXdqNFsvfAXVWtMRQwVnt1/5eW3pBlzxT/ReQ
tdVN628KtXOZmJM1hlyNw2TpV2RmT8yhUNbDgoP0wHQwx1oLzAeWa9cK1lRahxw/yj7KPKYkU1Jz
qC7q2HNBYZIm3e8np3AL6Ycxv1w35IuRJdzB0MWqZ0SWRAxYJ+Pdk0dL1rhlihknZWg0E2g+P5eB
CChC0PRr9XHGuP6ZuTxDE9Td19IqieJPzOSTsEmSoOqFo9y8Ykf/VjfBD20o6mFtlkArV/TFA9oK
eJm/M01ae7Lwbgritgkqk5aek5gNOQCFvyxIIJ7d/kTmhBq+v95NC4BKgplk4TfyF6A6MRaNsBu+
o+E/Hu4Oo6q0q5o96dEz85SmRKmEWNhbY0CApO0f7hTeTsU6ApnnjcuDrVCO6+M7TKiz3kEBVfou
YqmZAEz4yFdiqe59i2XpfMeMyyaNNdATrbNgnw1ARyWj2Ewy8BDlHTx6uzpfm9OA36y74nv2EgOT
Py64oXB5qVCdVOpiLQu0SHMHg1fj3n46y44JFBSwV8MuqShO07SAdHwqYQrQZ1JyFsyM0k+1dXer
WwPk6dtQ4vo766znxFDMnKXxgDbAbNIUaORm8G5ypor9lcvmcWBklrjCWcuVpxemtGfcyY6gBVqU
DPYkqAGxRxEawYR36oEGWgjwsIb7W0PfLEzzNA28xukJSraExce/q7Y/ZZnaUTo8227uEn25R64N
X/r48MB73HL2P/iEXo+vis0Xx/zKNUiFfUVP2lsRlEbkKSWrSIS2koL+sW4khE9X09+4Zgsl26Hy
wBCp5KEYzmfa9tKs8lVvQ4YSzpw/7bxd6nLq2Ea/jdfypNHqpi1qMAGdoi+QlQIwKO6WS8MhJICQ
YigqcQ6U7zziIklVV4S4VQXHMvcGvx0cUqYf9SUXqGztD7pUdgnka2DS+d3q4wDieUqlr6y9sr/U
7JSppPb3+i8eHAakncCGz3+YVd2VwHmarXW4ep2SRjRtAIhEzbRu+74+1SJnxW+7GUyebCHlgKv0
h2PqVTwr3LSi6nqQEhyC09CYMm8aVXHYE6LU4nRp6OHHiDtkPmMAqV732cdHRRMYt/QX3SX7/v1e
8wCWNrn3HrwuZxu4e35LQrf4/XKXVdbDohlcjuw0KGAblIqdozJ384mWRavlsfh0cbQcSmB6AsfN
zF/lcfU9uuKIwAhi6u2vsOJ5iRlMe10pVdW67t4gR26nBiLLT9mD1u96yMVXMs1lgpYCmwLnLBe8
MkcbDowbtw/sP202mE2OZBvoU443aCmoGyjgd6rQjr1Wz+2pZMxiGjHY1TyPsGY626h4HjsW7X3u
+E78tT+RaeZwbq4Lg5nW4ewEPL3frWMtwa6Jdf7gse0keWo8EgDEyLN4Eof0F7wJyHWe9wdtjx2e
G/hmm1Ner8FRzkT/nBdKOYg3uVrSaP3srSqQOdfpV92XzQ0a9vRtpYGk8LH/O2JJi1i9/bvoknnD
clCI8yYoOUClBoA1Wlc2TMcbKvz4MrrE93C6723up+KL2OB7w8mD9E98euwiJBkHEHhcRzPYtylx
uezbBXLtJLT2doog7K+UM4A5FbdgQOmtFADAm5anpS8sPIGitagYSGlnFb7/7F3zi+GDtNLzVM9n
1q7FTHXT7dN+I+TCXhPdOC9xipg1+i5HY8/7CLmoG3hRhBihmt9zzIFunuGyFCKjBsFut3w0AUNy
FnIY+uiuIEhoC252ps6xFS5/97nCkBLe/ul8RYkRmaimlTOBd0SXsh+F9vKaHYucEpTjwujqw4gD
JQQPP8dewj78mb8ELwJamxaad9rzIT+7Cz/cFqNuAQSyMuo5bivVbQ3frAdCbDuYpCacgVKJLf3/
9bHuw0w9XOQF1WVdzq8fcyMwZy24JSD9WJbjphY+gHQnXPQT5bXaHNAKaWobc+0OTxVcyUveJeii
ocLmjuCWGhM5De0MdlILHQTZwF+US/Msf25eK3ouwjk/QpK/BLlyNs/gI7cyu/EhwADIpQzxtBG/
wCAT282pSW5MZDvJdkkMnNDTWLhdLkb0uxE3r1lrsDbPyTcxH1lR8olenPCVbR25k61wJReO8thu
9AgmDO0aTAJvdKNQZ/jaUVfeIxJf8Re62aJhPFONecD5wy05lC5zHZRZ00QOQ7/SFnIWymo4QvT8
dby1Yd28+p8F7xElFMTWJ9Vh/J9AOmbafiSvrFVF5QFiLUMj6U8G95x0X3jF8XX9AZLoK0xv4lLY
XuskuEJV3S9JnuKz/LYK+pUSasKZJ2eoucFBhIr3Vxx1x3y2gjvAIPun3uFnpuNZP9FRxxkHd3Ti
RkpM20rLOhWvz6C3Zd+RHblRBj1eUyxvMgCKnnWvfJsxaR10dhw8zmXuHbuqMWOYBr0sTgLU42UA
qJDxnDXqja/hWkB5nLLmBeaQQtPnrlQuO8xDU2TKD2BMc1jW7n6mCGljP/0eszFyPnZzbXQCkATU
hBkg3uI85dDG4PjUzZZso010cMdfrzrkUJ5EofwTgOWdM1jj4Mx9juyPA+/1FBIQK6MeV45HJkdz
OUosgPqLswxylT4nXrXjfoQQzr9Du6ytNyHm4lJSaVOge3Pw51UBpYyXajQMxkYaxI6l68dboxUz
ozVDqo5DTQOqa9r5Q6jSVTv2mfb1zdDfSxDWosLyUX58dHbS8QRAsFE8iCrHCWKV9tCksVeigNXZ
E1XaP0RlW7DcAzS3XM+meCcgQHic9HSXTu9y4L5pJmAYI8n23GbPXPWYtl009YHmmnoHgAKOORvU
PBBdUHvdQ/c0qtwen+HeaWxyek47EinDlfIfLmUmnOgosDcxp7Z1P5bavGk6olUhXT2zbx2BP3No
HaeQXoC7NqFFziVoZokZSTr+v2He4XS/QpSvDsCq4I5MHqUB5Y0+T+1+TmQipsvnb3YgU0RhAKHm
SPVztZq0OuHdQZ20HHtmdWwvYdOW1dgpCdrJpuUB12pCholslSVXCu1KES9/aIEa8GCbtBNiYLOy
UCjehvYlmXHYC/xrzhhmuTYo16xILwzRXR5FuSLYhrQ73D2fYXx9tnKDQ3nswxCCy+9cZZEJh+FT
xVmsNauT8F7xm1CaN8OxHNUOsNx9Z3aiJbglHxtO1lg6hmvJAl1LauYpNxbJkbHvck7qBWkqgzmz
Egu1Dsgt5KSS2x8AsUeQK8GSlHhQLSgUOSXhNdSKS2BQ4ukyJ5s8frGtlA3V4tfVqj8Uj23FtLMR
eLWaehr4IK2zD/rNskYEGbMWEMjGWqkIAZWmAsXgIGIhc/32vVwY7lIKn0Xgw2o0reOP8lm/jAWp
r0sH/P/iWRZuuJcysy17UmghDefPscOADpw22/ZDUefhqW0PKAmTQo6G3NvGMZZ15Ce7pQkYHDjY
HfQ3Zz3gSf3D9PWSCUOMBJBqQRjhUAEkk/bVLrjh68sarjLQtvxgVpb7+KwjkqNq/6IcmOdYtRLr
Gpk/W+xsbvSRGBkrYVhdb9DQNajXaF6DP6aRW5IkCZgBA1M9BiZyc/zsLl8iUpVvn0pIttBNigpa
X3/ZPDV+a5/rdB0dIQM6+7kvzJWlfBJizbA+eHNHNKvTEcjvILIBbi0rt8TMh8zFphNQ05BlS55i
sgFrVLBR3srkKEM/KOLn3vCsLYEgTRPWVeKJFqnDZepttMS8NjvVxbbGyzf9QTefg0V/eUJ5IB6q
brI0/4wkGhuXectssp/eTY4PSW9/258DKQDt6Bj8O7rFkgNwl+e+/WiZISuJwYWfdvfD8PLM6ZfL
SV/cYz6OuKspObagQQXl8rWKzexxpP3fTdWZWp6PlWq1H3V9juc6PuBpv0bOYUjJJaTouQwNpEzw
Lu53+v8kch4i1FiNY+fOZuIt1evz1vffHv1Y0b98zhusjCfuehZWIE0jwfNKY0bQIZ9f+vz2B1Dg
yqbT781QlnRZz71OVUWGwBWklSo0C4FIgOKOrOVnOdvHdaVUQseXfOEgNAQ6nQxwZmNnnw9w/kCa
kzSenK5eailBiuZRjhcSHbWiae4QTrKYsCUnv6agUEqgb9RLuvIcvjfA9nH8oUvCCast+s4cWRCU
370H0G1S3H6UKxk5C7svKz3h6hEh+ZL1UmxOu+e4Ia76ixXVUhpiizSlWWAXfLzyoiz5AkDbTLVc
HnVBg41F42wGQVAXNRE4+zvhXj3f2aBusM8uf5B+kBGangUVzG24fA9L367fWh5JawUr44Awmk4B
xuwlc+KwZdh2YzJcX0RhITsjLzcTSYAXJRdfRplr/1QjbXcoQQtvN3qcCwVgvkystqdwG4vHfJyM
sUNwFr+sEwAM6N8POOOc3oW6dCAZrAwlP1ZDiGuRIOJ4oghB/lPiUKM7RbSlR7xmtlDlUZJwktjC
f2oBGfMGFfVVeRk+SHiqKTXLW/zPPPxsV45a1ZIWw+0/fB/Ftaf/eFbuuhkidkFdDYBNjxwxdjw3
ZpRthjTrsyC8s9S0/MJ2vPkQKosDLW7GEE46QMBjGilZHP7Farky6iquUcPrgOgRCnXo04Q/4qiK
ZbljWs/foz1FJCX+mBGO9Qmw/+Ad93+ux06a1fHlHgn1Np5Bo+rAS2aaxqtjmr/5Yxi62VBjiIp3
Jba+QrY2QlrP6QwTY3xX/4uC9mAtBkfanEWupWES59KK4vS9qoUO1b2rWvHgdiDLW8Yz4Qimmgp0
rZjZ7znCegYuDYMKt9OodoL55/r8m8lZampnqUkdFW4avDx9V1LjFWsse/y4Avwnc1i8P+7M7Opv
3DG76cIBeLd2izNqj4q7XRobTaDSvyg7b/XoEeNkTVMFOLBzRfN3+HgudTHB/BzbtuikMkn9/ZQ/
7Rk6hg878wkYwkJOuqEZtx5Z1pSfHmqVnW+IvgWnFd1G++zcKtn2dr6MqZ5i6kYy7RR45zc/KSQP
sH0B8Ao2NQam0cXSV3qn98uSzku7Xb2xZujaCgMJiH3bnnUQxDzL7Z66gVUulM/8CiXlUCUidifs
p73rFiaA0OZMyS4cV6jNFXtxjKTiHmOzYPSPkjL+cddipP82FYGzbLzqZD/UK6yAR15KYg+HVRG7
8b3jSbQXIRin51Va4Fy8eWrukLyaoskgfRBtmf2yGQazcEyciE0LW1EH9HnUZa6NPWfAJmh6OXTK
WUFrrtpIpImzPccrwERNLCa4MpbnLMIdug+2esrP9jOGQVYn7n6ozzWYaCRYE+YLMAPDPefreLg+
pJLw8mfVf/Y0ZBb5339WBhpJ+09TpA3K3kKrfRopaa7OBsGmVgfN0DuO3p93FuFCozHAPrm14Qza
ViE374FI7W0GzNC8Vp2xBVkdlHNfVJutIlJpA9eL+93SJlFSKWXzhdLZk0GdsT4FdLKbfAx0Gsnx
B3/ig5Dm3H7rOeR51iEdwyvszrx0pGF2sDJwRb0FTKUx+2lnhRm5jBi6CtShlymgALF3ALtujPd4
MNuHUHCcw8tQjeukK3lVixGTiBn+Hg50Us46C6EjunnFLhbFr8mLFePEZUL7tIJnySN6oM2IiyVM
zuwNFpzQabxC6fPNHtCodGz32v+Gu22aMjcZaItwq1q1H/Iwg2bwhYJVQlp7raMj+4lqR1eAGQ3j
L+WVjBEPT6xE1U/Bg3JgXButp5aeOfeGtQ8YqqyYencfjYEyeegcDJoxlBE0PY2HUKOJ00v4Rx5t
kCuVT65k2kdR/nEM6Eed/jb03cnw+Q2VVj8GQe3DNSyFJ53Kl23tpbWFVrGHMLOoMonl/DucndZR
0b6y6q74WvmsglgmdFvVlkXDRZH7V+5hRlYht1Kz9/1Ftv+q0Ts76Xj+Uvq6OIOaN7r7O62LZZwf
bmYH29S58koHctY9jMdauw8n8QVxK+y8I4acpQcefKz7qTuAyJR29kfD8Dk9RurrhkbdCljipAMs
by1Jglz/7K2BGMHantSon6iyNSitnoXOPHAY4KjcsQc9l0kQd3+4EJL08dXeNA+jwiHvjWqNClw1
dZlS0Aik3ls+t76Ib4TAUmu2Nv1IDjXZadx2703Vn9LXNOA3OpwQYOidgJ78haAXOBO5qPFoUVbm
Ve3kw9qQdUOGnP6H9LhPZm1GCFBTURtUDlWZbrjkJQ9DbaaQo4wKPTD6ypkY9vRC8dqzZ8zvNQ9W
vaa8jONWy/Of4Py6wqemsfb/E6wJRjrd+Xf0aSlKtDpLi2pSSZ9D2zIeRYqCkWCmSrBV23gbkVzu
6V/57Rb19EG4nGEwwNqAIUeUWWn4493OWdfQ3ZlK5LdWrZHBCV1rIY4RJRalB46aZYk/hsEtA/eu
5JAHMMFLEPUg5JpWAzN1ziM4+kWTz45W05aXK/e+G39SkMpg+by7/Y8qiWvosoNBVH6MK90/XQCD
Lk08NcNEbV+nc9lYfDb9lRSLZ2tOYtV1RDFhhiATZ9HhRdQuts6pm4PBeXirSvjSALBezBZMyTB4
ooaSGcK+trRNiIv06nd5yzOslUKVXHOsCNRAlzA9wEPkSSQ7wrNkVAjSQ+l4lRDiXrcvyLo87s/8
UDMadW5yY5W+HBiScyfNFavEG+kT25Eg+QuYYrHUz1ifrLj8XXCNE7e4ajeMyC9QdJGGIieyhTbS
oOAe/Sd4RcxpDQkOj/Vpt5i6efku+sGSWqDiFVrgmWBmiSaulnWunBDFTnJ91FhiHsJooL+pa2xM
C75MehYrZ/xZcW4eaTzrAl8r+hhlsIQIfNLZeiipo4Ki7eVpTrnQDKKaxtuudJ8syaaw9eNUaBjR
/6aT6xQ/0FsctQMBul54gtqFkPvyaEiP43eaYPUlV7QYVY0+nN3sbVW9f9x1I+p57V0yzdalidZ7
nQ8IXq68zTK0PliRZ64IKosn7d0qOq48RmgjM82ls9MyER7f/KeIltJ1z9iKk/iAUmliTf1g0X3/
dT5L9mkaLQfU18x5IAn5aiSl+T8GtDkQEeHPGBYE1Tj73cS6GRSMhLsKUnj5CknFW/1mAduVq/lk
zB3vsCTVrGJGbpQyiaWsVxn+4eUa6LCcexhXDAz+3fBuA8IjC0MaZHph3m19g2PZVCx2FI2F02bc
9kySTTSNovNRBZJuVx17oD3YEkKMdonBqkqyyWvNOauU+WWsvzjkXO+dQjZVCyEMenR8H+MAZFsc
VYkkgSNEKBqLP73nIFXbp2uT65j2E6x5Mu8xH4w1mYAdn6QvUN78E4rDmMnDA0gIJANC1VUXo2TF
te+mA0jxcEQbPLmHgKpoEr7Xz2BSHJhUtUd4hrLTQsaauKSnnitiYMv12/0On/4ozSv77rhYvNUd
Nqpv6zXI7MHTuWXUZO63S7/m3cnUu0tertb/4f5rgDClStqpJaxTSpquDgA+bpNiLz2b5X8ABPff
jfxRtY9hB08W5LzGYSFPcn1vqow/8QopXMpXnzXDE0eZ2XsLAjuCRw2RjHwpBghdMYcXFgw4k7q+
CpEi6SEgSUaNuQYz8ZIrXdmrUBDtCddkE241R2QgVVKcPfAr0diCBi6unmY4v37cIBpzWTg5aG1b
D+3QqQiBOMFb1OoTwmVf2s4li3201OITxbagqVPj2Bh+L6Bz96UbYFebdv4JovyBFsqmeyybJgsH
3dKrnHCptbT5NR5L3I1pw80ACqfJ9H5JmQ6/S5nSdNOFh2ojw/pcS0gqqJtysg0+/hnG1n028l+a
6YPjN3bR/Jkzo+xfqpvK+L40RpTrGqroTSylvUgm8Rg4EGLnzMONz5WXSkIxM1Nr9kf2fNCqRJw8
XuiT/pQJEwJFnHsSjurLR3AJNN83QAW6tLN3Xf2I4Be8SFyRs8qskkh/U/y+B61rvQfUygppIe/Z
yV63I0VfryynmuAASmzkdP53cSblw+7RcvpzM02wk2S1h7uu1Hhdx4yGCONpBY/fGyOc0Rjv8BZQ
ZAf0zqnvNm8tjrErQixj5RDS2erlmggmBlTYyqNjROy+Ahv9WZtCU+w/kiqjMFlM1fGwS6k4bE4x
Arx/agBvFkogD0FuSNUpDI1QWWX8tgZcxQqDjrx42RkrDKjAlRbohUMENVGF9RgA9FxqocDLTXhO
qZEtLJCPv3s0tDx3BB2N97TMUkjUIiu3Yp2ZkRMjKhiOgzYHcBNbxK/YB8OnLRmQs7wJ4+vzDmM6
zaDpQlh1KtqHPBlYuc4m1nB6gpqiYY71GwztvFt+BbucMSVcXzTcGCJ3bxZCIM8+OcZu/Qjy0Hfl
b8PLmCSu8H7h52zY2qv5DTWrQoJOly3HAMP3TCXHWc5cNigv2bHBCLIEap4WWb9gxcaPsDxyL+i8
ftfcfy2qiA984mmCQMokmKUYi4lwHMAMdj3y9F089stq93gmS65nPC8G1olIVW4Znqta/kgY3SJ6
vsJz7qQJuVAiYiLDN4f8wIESmIyy9NdSQnJ1FJMHvfiXscMSMyvu6fK6RIXlVg5S/FNr1z5NJFjb
M1tvFg4I43FeqEywjp3TYbFMKRq0qYpUhfoJpPnLKcxVc0urW172TqpzGedyrsr1IcAD5zd2kTA1
JATX3Kzs9/Fc8DST73cJUZUUyEY/s0mjTsPp0VfYLOHQEtsh3s6l2IWK7wHXTPy0QaBDj6ruZsT9
ZmqZYeEbAipKG57eluEtitrCoS2lAjmf9OARRo+muaPCoP4lfeHzup+RBhtNfyZQ5gnNEpT7Y3XQ
YrWiTaP7faiHTHyCwQAAfWxqa124KRFwA203qFKyseWLs/gcfISImI5+8vzuhiK+lms5NIoinwCH
SxkloH9auwD8FCUXMFbZnAEFwMx0IFamgtIZt2Ha1BrqUoye6iLRBRnPvHTyWfMTAxB6flGjCLfz
HVNyqSjnaDTKjmD/IJLDB8UZ3eDcuZgJ1zN3/JpC0E+0GT9UMxgsiwlFwd7HQ7quu7c1heonGmse
EAX823+OumIQSam4toL9ryZoDPydkjHWSo8J4GIyQcKem+EuRjyD3qRRM+2F/D2rwinF1CpmSdO2
SD2HFp08jyovy2tWQr8EF7zUDSgQVCKQtGgbxQFXydgE3p19fzVtr+DsagGPY+9NrVdIpJoX4HLi
ChSCnvub3sSJjpgBeiR7+AQEUghv7wBBFFnA7rRMyN0magVWNkOuW5sfd4UHH4foQg4a0W4WndAX
ShVQPrFKeez+SclP2Bgql4yQl6TFAuUlYgzfcqZ9hCRi/qJHAvg0CxNpM1MSt0LX7c8pzuJCYG0z
LR3kfJB16F4yls26n4aSIcqKdnCFVibo4yD88U+7YDvV3PEhnplgPxxKR0JDtao/pbJDeEb98Iwi
cTMDfrhoA9tVXyjCsAqRM9pBmhvtfigGnxIB+uhTqx4FNFUF9i8K0vgXwT/qu9/9cZ9/7TB7NgeI
O3wmX1FDo1+vqlDviB+mmMnuzdI1NAAnuVdU7q/goqSLuWjgPu0nCYb6c5ILnCq32LlxCtN6xexy
9GfmralCkgvyFazRB2kNw5OlSy2FUFrJ9nHGeO5qZQu/NRlsj4cvOp1bw3EfMiKKNPAwOlbzFBcS
4PC6vCbNDLjoKwHZFeRn/im4tcmvsx0LFlkntHEu+R0brRvmg/6qPUWE6qxINLSBZ4OZy6fSLiwH
9hhWTJKoBpSegZ5K266y+zH9+zmrrEG4uvDOcBAn+s9xk5GVVOGW+85FF3NajB1nWN8FlOfD/YB8
YFqnDMvOp+9bAB1nDer4HUvZBfF3d/1m7DS3wnjYOv6RMcgqI3XJpoa0lJNMm3X+6kQyHkfvaRIK
izC/TwOqcEp1CXoCQ67pCDrXxOWvNQZyUcI+UPAqZDop8pwhe9KqE7yIiN/UChM88JQbwt9tETOx
JT1R9MYQv2N7/5mQiBaks3cjPJbo1Ewg+9v/MTpHltJFD7cGJmrR516uuNuRgam+hWJpOFyCBJRP
htKvm22paOr7l7KBM9g/WgJ8V+dLY6CGGhJVjCLri8y8QgYqiJEJjRgoUQ02sNYCWKdXlLU46L+i
pK2TXSraWT4anGNumooq0jLY3YP+haiiv+YtdJaDZdvnaeC8xB0Nzbapps01MIZ6rkjwN8QffcSp
ZfJcihrw9/3/EzrMZdllyrzLxpLmIWP7Z2LXZZFbL8cbcgoStJzx/0tz/cfzGy7qpQJyiC3oqRDh
kyKLycvrl2m1mRrK5G/Zpr7kSbctf7RH+cj8byK6mhe4ioEvbB7Llp+keTulj7HE3bIGPfm3v0C4
oBOvp7VAl8YdvebjqDVXilE6sLq2KZe1nt9MwH60V1GRkqL27TVI0LBvZIc1GqoKMhS52bZ+nFLr
JAskYVNZXsLqRWPp4i6NYbRIgrd7tJO/wmsO9K7JiMU5axUQf9Wm0fnMtTjinZj8ePrq8OckZwE1
equNNo2UBS6Ywi+9EEg2JfZgPaUg8yskm45LhjzZ5ptxDxu3DdU2WRJmbmeGqf17Vr1+jIfGEjDE
R/YzDx8/P7oNeALfCYQS+h74uPVYI8G9or3kQ4RtPJ878zI2Q1QNMyRyGRzGam5IGzI+yWAHoN/i
pU2/5/qXQ4Pnjcko4YEim0fbE+Ih4guvepm2BBBLy30kJqX3YjUE9AJR8lY1NO7f4Ou+ttQ/tshs
BiXEgpeILO2YxsYTU5w0z2zw5kjidaLrpvCh0MvM29sBk9Ul3sdi8moDKMJPlXEBA/xaPWDJ+1TG
zTkk6CivLB8ziyUo+SEpC+fdg57ZlIvk0KlJEVtU08sFiykqFRpt8NEKsAeEqMczlWPFGVq855ce
24ghFvcrp2Ed1ppiXKAmw9j4h98NrMqX4LQxzYEoo5VdE5HUabsiK/PYUcLoZPrxKPYcDA92QtD7
ztRGnw87gFofI+IPHvWg01L8LO5qNYgF8+w5g/HVJZhPS3s5GoaUwyzwbr/EOoQIhSUNb2xsm9QW
wIFAitE4bywg+uZsuqnm/DF0FPxZ+N/UjoKF9qEr6NNdmmDKp7X3A1L6GB/3sFq+Ce56a8OVIPJO
Rq9uVbeo63UTMZv0Cp8ilYO9fbnx46kKjpCDufBYyeLCBwyTL5nPHhgXjVkbM+I43smXjqfrh0qt
eMwHLCZlowRpeWi/2jEuePJnNVZov53B0wDHGvTz3k8Xz218mNWSN/cOJxJTTPvO5zNJbWVCIClK
+zc+5soSawfL8+akNdYXHUsIA511kgGl/WYoH7rahbSZTlRTlb5G6PbSM8NqOgnNZisSVil8sj2n
2Llg0y0GLSdujTxiSjbOiOVglXkkS4muYagA2f7pnm6McKtHvDCbHlFNDTfUajGvZi2+/saUD5tt
3ovW3TabdvdtZxe4thB6bSd6NpyYj6R86aoAsp34BFrBxtW54Q+/sAs0ZRdA/fsloehMZKmQ9LSS
27rtE8jztc2Ri0XdvLdNe2EWLSEp4mamSb2ZXsjP85tIeb6vKnXR1T0a/iYRQrn3tbaXfvJiMVBY
QbL92RnLXJk6hayuPFkJQhP5VBkCiDtCC7K0JM0ZqSgZ4uACpBYdgZsLd44A/0uGl159cBIw/rjQ
MHWHp8wt3UiloY5Nt6maBOk/nwLwsGAMmqsbw8+NxF0fvaumwYaE+kQjLP+KFmYoqb2ugAuS2QsW
aInTVKUnwQZA52fgjRIJzpmdMDd8C5goi8WJPIWDfQS59MjEty+kTGLeOYD57QDjL1I3MDkxAaDl
ZfGOrOTasXb6eXIDC0hR3EUFeThJ9y5lROXCzOLyt87JIOeeVarQGovTpN9D3ahCmOZKfXiWp7KH
pO4Ngk3ZlvnttZCecIhcjx6f4X6mVTqxBKHhciLF+BP3BBwZ9kBuN03+O3jx8Ef/Aw66PTj/WwG+
rIK0FnvnE2V/MaBeCpfBx9KZ9p+ofdU+j+Yo+7FyyiOrB2c8gwDvfOHn1RYIviOZbisK0pxFGttB
+gWucZsAq75ERqJCaCW5num+wJ/Z846Eno1MSKUXS3Wr/42H9fdQv1NKOTV6ei2Kq55ns3NX9MkN
p9j4A0GZIWJ4y4o86Gazd8iBEE3/c4VYNnHr8ixWxUkQBKk+yAgH2tj/hlIEcJiJ0thv0MwTvxNg
YSAF8rov2FEL+jNS7eTZax3RINYW+ITKDLBJJPELUr4gS0GBn4nXRoLD0SZja/80hBqXy/th98fo
YatP76b+lX34WjJqMX9PxGZ2qX0muQdrGBW+wXfHMkbxcODR+WE8ItE4lI6eTuX+yNtOksEBkcwV
NPzLLRRHcUzxelLnuBvoWa74Vu4FOpNeudnqRXgNPN7gdW7ooCD48paojMLwbse+zubb+AAEc0SX
A/ojEYeNAWWPUxQnZaRv7dkbHh95oOIinVbhT2FbVKkWUCbGUKO91znK3o77BK7Sa80CXPgZLrM7
OdTIW3Jp7y/DLGAsDAt/HbZ3njc16ogcGLNwiNJm/1fxJ4925zvOp0je4SCSpzC5zHqSG5CHPtRF
aAOCEvkyoUfMx48p2yVyU3sC5KPsuQa3jYtp+9XClOjz4a99q0cD0dnI1P4iL/bozL2pF2qgYbJd
N5b2o7zEdEFXHOQHOfe6Atcsyr3pCqyriXHJ8ayZN5IqW1XYrT3Hg5wzWM4NUnAoj30sO8vYj+pX
JVGy9s99rKcbUI773Z2D7wNYFCuZrOuQihvbt35t5uB4ysUE4tK7/f7Rbd5o9x64Cg8uGW6ydrT7
542/SwE+n6+Fs4u6DHG4dCWTuH20B485MFA5RZ3sC6cCzXu8JBVOXqEKnDx2Ke5v8/4YiJvzxZOq
7oIF9HRLWxXc5VYKLKMQuTYJHON8RKYyfJCH4A7Rv2Tzmx/MsKOhbZqql87w1jcZWDSrGtpjewo6
65kmQRFrQRDbeMHO1mnwSe5eYakGP1iWUgKZnRT/ivwOxITx0j5BEx0KlVKA7qVMK1d/P4v3r2Nj
TVxv/wuv0V30CGTtwoc/DAe1T7jKLiKmwZ1euWTw44Z1RnWyzdcXz5JtLswkpYhn5EkYFjhEkW2U
WHlDL2PZcqRcJlzMtFw1c8+mKYYJ8mxSVN5olCRd1yqjTsBT2WIkyBucw3f6zGvVCmifMRvTNaJR
EU+ezhBJEYtwkgTEEk8RM8iE6fEKZvBmk1Qr5gZ4acqjRLyEoIdjgjG4IEmjFFgia8WGneT5UF5H
O1TFg3WgeeGsMT1rgrJTVz2JygyCesB7bu+veGt40dy6IS5A0HfJCk7yKeZuG5arSyx2rcf4Xpcd
1BPTZSYJo6lm5HnWwR430xXrn0TNLc2DEmEtvnpLs4pM1n+/vNeTvKs6tsCqOz9PehzI+ChLAk+H
1iy/t3SBzYHtkG6XiluLURVUkkCfryFHFJt5ixs2eo7aph/ltWRnb9sBodJnVpmU5H20Gf3u9Q3L
TYjRbYPv1+RdKXc+h9KJC4EIk+1ctHqbJqnxdiICQsRssZPnz1dM2nOfqBjBQQsQRIzUobbjUpm/
Ch5bE/+omWdR2wZek2zyUjc/4JD13GS0wAD7sd2i5pRFhrugHmOaJn/dbsKkbd0MlZ16zeyCqA/i
p94s804IRSlFswx4Lq8s/PiY0Nm97LsM7w1ua015tKoli+DPe9R8xeqdqYLw7bgYcdJZc56VzAPv
1kMS+wOoSCTXrc30TbJrJN+VYj3I5XQWUQ15CYvV17MsM9tnMUfyXI0Hhe4FJelRZ9yRXSjmKzA4
3BOM02Aj5brQ7yqSnyrgKvVfnLpUGlpYmsf61kHg2MFf68JHV5sQs6uqFsJ9g/MnDCRItZ/43oNe
R7oNikgLT/KTr+7IqLm2y+ztQ17e3QTKuR+v6nliN0xwY1XEcgtZ0FZrLmvPVlGbMNsBejl14WU7
ndeXa8/romOBozll29an6pqn7Z4NJrPP7tF/tlIhH85+f1dpoYoSZHTuFtZ3EgQayJ5izlLcTZIL
+ddrXuU70+mOgybVCqZGY7kim1STJWnTzM7/k4fEBOgm4i7OnwQhlihDvmtRQA/IIMsjBaPp3G2V
Q3UE2IRF2ergf8D0/tOvVJ4YzW/y1mnww/nFdDyPsvYuMKdRLi+i2az/JCHpXpE0txyyWnL2GOhO
QznPQhjRKYLIIByIDHpJQEUh8joGtSIWsQ/hvkG/MLz5AfGRj+2OF+KhWMY5AeSaLw7ItBsyjEKs
CTlWMbhaNFXISwE+XMzdSnAK0uthn+7IsuvgEXwFqUEebHA+YZFjY1PYuKE/TYcLqMze0THSEdPz
LQvvNNoWv7CogQZrOnxvtOeDP4EfSYuEZVrOpD3KaZ05cFF4eDcvvZw1zOEZe7hMuOx/lZq+VIX3
IQkuDMUc9vstI5ja06na052+q1WKO1O0i5MSSIlforuFEfCkzcNhA5co3yeYjg4xTzWZON/4k+hI
ZRMI0UCex0w0fwOzl/vMEuZXOJmnqL5N0x2jLG0PqXBAZAdzmJe26WKzvO188FQ2rQ6ekJv+3Ahh
gWuxSPXgLhDrjMK3NaQAOz7YKEQMLQ9zUSoAAiPCZ0ebhdOTxIytwNSBvwsZk2sqgure3xRVm1wn
1/hYtyPI9LCLlcR1S4wGHVw55iteHL3+iSveoxgtrVIE9OMwRbwwtCLajMmNLkd97pxX17Y+QqDf
y1GDQ1TjNNeqO+fCJAuwriFN0TiQXxxonNoQCnUpMcAaF0N3qTnVN9bGgBQoSd4U3/PiQyGZ8WHg
+5v9UhnofoNg2BnYs0Kl/qMV83QDWXHdxr2Iq7BTjaLAoW121yOaQpS3YxmSpsr2hCtDOb9X+5TG
GH7Gndklb7gc0bgnEsopCytfaDlXRfNuvuYwTiJBvRjZ+/Ha64LGA084G2QMuwXgRH3FT5mWXpky
kBan9f55acDB2M+fBK+agx7/Qqi51hyP1ZdrJrWTeLW2WPk9GdwtE70SbycB97S0KtUIbiskjWNy
vqztw2CFCjfJNNKTKXbQ+6GwYQN/4dmMImXQuOgfJRHJ8Q9t3lKyvqfOGm0cARAKaMfug47xtIuc
oUpFrz74pveyMNUtnpzbtmx/x9YQaI0LEHBbzi53LWr1FWEltAfnwp0UUBR6qfDO58u/8T31OT+L
nTwsq2z9EqcHHVRwtit2BBRXUPWtdN6JeQ8BDq74Ht3rqihqy6wC3pcoExwfXcE1WQhDqqnoPJjn
kzq7zuJOJx6nm9hUbVTRoSmA/p1ybXeakj4KfKdp84IAKMJehrh1Ewmn0d6H2KkIE/HzwpvK3bv8
IVqSvVCVnfDekciSA1Ms1hRjvGdmla9/m2oJlEbC7gtbuIw3vjrUgav9gD/2WqX9vMIVDnojqhl0
bqz9yKJYembGDW2RpeujyITrMh8XfIrPeTvni2Q+aM9JYYE6iJqVG4cEe5/sV0TThqf2G/xQ/0q0
1B78a6xOfWZPTDbS+3sop/Q1d57c8GM9odejHMtnLmVUftIzKUZj485omDtihO8pyecnCspL5ACe
BnKTpFjlmYvXAIwE+mzEGkOtQFGIlFPl39gfFNEbYNQO8OZaySevuwyA6jaSiHiCQjWxYQEMdpPM
GMy1B0EYVUd3XvH1+cs8jw2RToSAmwrG7sJBgqfWrFlknJhK4O/8EsifiXVyaK16mKNy60omwndj
310OZyosgpjHixLc9lbnby84gN+JZOtdiG3p+dAVMbrX4MysJIAA8yyGJ8C+0e+zfytgsQurDjBZ
cWno+3lmtM1I437xgVMxIN2vKexjKu5b1dHW2bl4hTaBHmG4h+0XecLPPsW+CxbZXIScILhs+gHo
aO5rD7TpbZ5KKwgM/Ocq7yQPwSHMII7zWkdsAeImhonH2QBLBa0pAPPNLQOcfgVaRa+xk5KVsUXC
36WAeDoM95H0Am3bTx31Y8hg9bqCzyBYW3Yqyxqau6v+avbCcB2dTLHRsH52DsZb0JDUWOIgd6Km
6O4QtNtv6q24VJDICBrAdqeFbAHBDtyyyqZhwEuJr/G3pneH6OukaYzc53069Sdtqu9O3xGTYPs4
yLk5YToP5X0Q8U8VzaQSJzG1ifesxfpfI/dW83SQ3vVA8RTot6Vemza/3xdSWtGaFnmcGujqbFGn
ojnwbPua8FIEVzeb8GpQO1WGjppiyjDi0GZr1luwnFuDJY6JA4x8kEeMKjNZ7LkV25j/t5xYlEkv
TV4xJvybRqrkZkXnK4mJbqTMLwtoXy4zm9gtppNUYdyL9/A32FkErIfZvaewVHe78bAJwvR40KJo
1yEPnmYkEkgxBGh4vDY8MHIpNajKdb0vHnLbetkzZmBY2TiV9JmLbWsuwLrmnDlRmLMj0H6uBy8e
IjR6aA7ZmfOr+xv+KAgq6phOIq0SJQ+EfV0Y92t7F5MQL+jLEqH5x52zMZtW9+0gSXuwpOHTcEcV
Z9R1mFa/GhXgMD+m8sMGpIt/DaHiyRYrkQLYNX+Q5wojeJEuE0YxL9C4VcILxAxWkX+rKrwRbPDz
vIaq62NntaYVIm2agbOW9nEyqPy+uFg12+8lo34OIdSU3snbFDeiBr2UfacNyvuvkHAbtAG+T16D
8gXj+V+rKtJCIqOVFkVcujEDAzEqdhxgEGHz3SH+WIhXKpY26VaBtHTn86l/xIiiWHF+5dk3ioZm
pZ+tNRSYiKMZ0TAVwm21rws8Zm5wun7yqK57Ui7jXo1aZB9DyTHle366QRFs+h3mwJCy0pkk2/2E
0e+BY0YUoUJp2ACQ/ENwMHSN4AXmC6ZZcQudH8AZ5hzQLG04FtQhDt669XFZlIsZcwRW3XBOBVLM
zBzNCKAzDWnd3onTj2/hh9+qrQw6U8pZpsPa7HFcaYru3exsCaTOAN0n+MYOp/sYi52Sc/K2tenM
VlF7SiZ1hwewQ7UzMF4k7hlMkurHMnJd9I51C7R2xc+pE5JMEQRRp22SPMaXmXt43T+0jVQp/H++
xMRPhy+izC03hAygfPHbOaF3wfkqwMpIjiMHgZTJ8GLLRrSQ3aiUfhPOQa97V1IvKK/uWeIZIlvE
0ZwxkhigiIGQb6sSgEBgVvduwGDsbbwFhTxfo8tUfCqA254FirRoP9vjig0NdUGbOih8PXBokKwz
sWb4E+uC2wsb0bHJ8ngaVcN5wDSdhDwyABa99Q/+M4FGpXaXG04rUsx8l4yWOJ3F7HJ9/qUJIP3w
UEp7nuZNjje4jumYAG7HkX2YvbrCrp8ng9+OpvBAPatU7QDxFcnGtN4UmW7pv828sCBtU/Jnn73U
+xQtx9tqTOwgUUh1NwWDPCNfs6Htsz7kTW8E6jxT9OiY5d9dRFGY/bj0AR1T6tgwGSniHFmLeJjX
ZfEP87bFk29OPTKi1szcMFgfA8B5UMQE1Bm+7Lms2UEUXwrgb2tksPltD5AKiQeTLKUDjeAdLHex
Z5bAmlrY0PqqsHBUAn3y/w/QhEggD1BlBMtitbXc3YFPcdtwxNVtg5/v2Ju/JlKwxHZhNT+rFqya
QI1yOC3+uDle8qAOwRF4bYBOLWV7OQV9IdGLTTX9WqOEl9jK8T/nqpgthxCKjgn21vUa53BmxplE
CiHOCytYUVOQwpko73chwuJNAjN8zHtGPP0ha830IVoc7qj7i6Y/niceJKr1O/VTeU+m1HCCqrTG
77WBncKjMyVfai3AW5MsayGC5EmyPUDb5/7rFDSZ3KsYLVd/bT+sylCmNJT8mg35+n4f1y6kYbsd
T2MGR30dvpePiEmy36S6ZebYy6mEaL0BGdZ7D+58BsSIx6ILCLVACxg0COlLAwHm0a16VzFIPth0
qrZEPGqGQMPbJnGUT6j5BUM7MH+MyQfU587rWpHKq/o976KwDY7FliLI1/IVvOwtf5VULA88mo0T
SZ8tw67SD/euHfJhmDl6J+RvZT4lp54syHByyVw6pLAfnG7G2ZalpHAUZCa9VHoBhs/YMTmYRrl8
uNNsqJoeUc5fh8gOzEcZtblTw8L+GpS3QZkCycz6LOU6jCb2nr5+TKOLMp7H8eXDXU/RayQJLOYa
FjLndzISKrlQG1OdkKCeSp7yzl6RgtHuhjRyxbhTt+Vd3MTzGTJVRtY7DKuT0LSJoMS+Q5nyFtJC
cdsgNIytWu3KgEQmzPJN1Osb+e52+c/NjAwXAPezEWEVXai/aGoRB3rslauNZTIlITlnEWlo55hc
CwFnQWRV0dtdrUljLYlnpxjX3aGlm2CEOOfJ4RbTdNtrT2UxRGI+ebMFsWJ5ks2a2Atu1qQ/Sagq
gE8/4wRvfInM3YpyWzkAkfXYn5Im3M00iBFLDWUEN3pfM6XpSkzLCV0NJEWzN4eWLYFU6irM58s3
gJfV3e6vmv8Iz8I41ZoWN3M/95SufkB3uf1Zc1KZop6u6Ln5pN8XJvBNyPoX+7AlkAHAXqS93C64
ooV4AhBFyAy3LS7LXJ3ow8vlcSKt9kk1yF6nSeODGbaMSHwYEWn1zBJAz4uT1NclynSBZJznakeN
dZicSrxSI9qTql1kurDM/9zVqgFUT0l/5M2Qfix2DdgwbnwTlHglrAaMMkN4mYmosBy11EMyL9Gn
yZ9uI+/MryO5un6q4SNvmb5h6yI2I4YmeinKAl4bbobQVsXZQBwgKuJ6Kn2WH5xElmiqdlpnu1iZ
Bl7A3mLRT4dLU1fsBESOflW+00DjuRCB6TDkNHUApcuu0IKo1V9QnfwEjiKrgJ60AsTkImMABIQu
OHOB6I4R/uMS1fTEtHO6u2B1x4GIZnuXraFT2Ee0afmy6iY+FvTaUS2Jk2C97Nx8BWpmICYOfZF7
mbbahbPhR10DmUm3sJKwcMuqvY4/JPG6pPoefiZUYhyzRGNapqNlZCgLDYEhV8+kYbeN6ZSCxjtw
1g31Lkx5blYvuuaE4e+UU6j2d96iVUvigufks0OUk9cbezAdZl6+n1KbBHA52m8siIRRJJ0kfaxg
xw5oGwbNy+Al61RRwKkJbrCXqc7HtBO6LmXEevERc0s/2elcp0vfqZPzTjN3+ysPFVpqWWpU/HYH
LvsXScr66KMI4zyjGcma7tZ1m1gVyeUP4Do5eQATxFTKJub/puxH76pNdHecZ+zJxxp3MZJwClzc
lkI1aNRvWcGLzavF75iXdN1BQ+AgSSSJ2bqT4hckPwITQUoEk83raOIM4XyvwOFvFNgejn9Ov6Xk
BBHpoxZFAnIYb3ft8ns/eVKvxszZxsoBL5I5eBkK0/p9FC0MUEc3Xx4jAHcfEapXWkeqyYHeorgX
+TU+rrNGTRKa9lleTiyy4X0ivkYFMSb/Q8/fZfo14h6DmVIawmZAbOfxYDji73D6aB/xnrEqmGUB
deQWJnSbWkOY7MrjbJGbAMTLcbFf54wjDOzA9Sy6WCsuRw06Qv3PLsk3qhsah5FizSv/Scc0KcmC
mcxVcZn3iAdIJDGHs6lwYnK6kfeYz1l0v98hvPdB+mSgow9xs13cyoJaSY7M5zwuQOwwYnCbxGDz
xUvYXQ/oCAucDVszxOoiW3+xlt0rbuVXAry2N8p4vNobxSUMm+CVoeOwg67Ww+TpZLKnp++6tWWB
5zvKMZ2oSvCkvNaNtym5eNV5ZCcc+tgqAb6g4pugCGx95o7NitMhE0G831SeaZc3Si1UUXrZWcgX
e+US5smjAoXDgg9cXzXZ3ARwJL7BHSP3tdHAHMZvhMv+cZSKqIwdOutOsE3DwswHpDq4vUX1qY2U
R6L3eY6x36rqQgOOu/VkK4jd9Ft47wnCQT7zZ/Ras8bR07IyLmlMCB/LEWoIK+EL/lu/c/sbA5el
Cc+HNllwF7CZhS9Oj1gsmiPOmE1+pVqQ3tSylvwMS4bgJPnVa0ND+rVK+SIZ+/jBRzvk8HOidvGm
0LzTRaW307VLGCbkpa8kkNnUXAqdruYv9nyP2cezuWzZPLnwKyTPt2oPL1rcDEg8bVDzv2sIRiwT
xpkBQ4OO0hIiUpxGfwWqzmkFK52+YZMo1ukP/kgPaPKlYpqBY0Fg+/UGl7ANr8RyPOZcRKNrCTnM
s+3LLn6ThIfbfwmVKZIfy1CzTxP8U0OWRrpnX4WQqljMg+BEp3cN00Cx7A2uXCT3cBm39UhzM8KE
tNmAGIqaCjUuv8T8eJe5FrtLHNSO8R/0DhUm9LyUG85vEn36yQgGVzkGWZyDzBUfwlOd16CKcspU
eIUcUQ4IuAoiexzH8gCCyz44Ft2kt+tXJ/yr+BtsFHlzmiC4RMEX2jTLQfEEjbgXfDsQHN6a4lfN
IQ4VY6jmoCQ18YYns5fe4FJ3tEoBu5v26qPvzMADqw9g/MbdiIh4b6RitVeyEI8chZ9DiHEnzVGt
/shfgVoEkh9EO5fW7FxTdWqRJo5ByqD0d/aq2qDMTIBxQq6i5OvIA02YJKux6EWY8fHQI/KwzLYA
YVsaxRLShrlcLpgCmOByN7tQIcFUYBtjAk/fLJH5ZIyCkTnIzcoDDFV+OI1CihjLHAMVsUg+a/b6
LTNu/JG1MIX6joJ3dJXdEtSbRcpanlsh5tI0h4+PSe3s5mo7sjko6/ng2CRdSO7Q5GneplPDLR2G
R5nJT2vP06Inix1DbTHOuq6H+kJPoi0DX2qHTWuXUq8214iNusNG868pVuSMDneYAAjn5SpG1jxb
PVeRM7deEtE8U2vNc1KRpYD7H+9EOi+TxN1Wi/dowVe6taSetknYCybh7/zE8ztMbGqLgEXRGG5n
wqpBfhQ3akX1ilMFSvVce7PCvOl1qAGpe7v3OeiaxbLblGdS6pyDOpwZWGQdns1g7YYYFIuUw+4E
Q8J0cpE1+w/fvSsDWs/OGwrPgDkZEyfMQDSvnCRRodimt9szXmOD4Hx67a8xjv/Zy7ym2w5FgfuA
bg6z0vjdpMO03zWBGKeLAqrd5DGuXnjes1KEt4UG0q47EPZBI6fARV26uo8I/bvQRpndA7gV4Bbo
XFi30hG1pQAwAQhq83ndLmvfqrz+WSlSHdzMh47uCa81JZpPd0APrA/oXYcOpW2OcwM49nWJFI01
klUol/LKhQDxhEme3I2ZhYSvmoTxUwY4EIaOWKhYip7tji/pBRrE+IfMfH+RWNvE2fHIEh88HI2H
IRm5R18o+4g2y3C04hPC8Q4a0+SGFdeHDmahsZuw5lpjQwl3sFPD0rAuA+jJ6HJA2WBXUfjxbBME
fYS3k8bqcqNk8h8U0krnrz2bCGKzmcxeLkRDFsKyEQ5shY2BVc4istPvdgDRgcIVuBWCyrNeFYlo
KmHWkW+p7GVjVsvNYQrXYNZWHdGyJPOBwl4Zm/UvWiWxjax3V6gw7hI3m+cqsYhUin8susGmwAhF
KX4qErRerYnBVvJAQUt9ecdgPbXO/uuWdu1gJir1doJJT+ToTav8xV1qduASoSkcFdVUGL5NU7P0
bj/5USTuU+NYy0+cMR0Ome1aHUWcO9ZinPjQVT+uMd4B6CKY2K8NcXnaUOYdb6eL/OPz5UHLqzfg
GBuQvcvlPlN+vno34ADUH/06/T4ssaiUPpyrrnqHsFzsy7fgIr6V7Zj1pe4cExIfatmy8lbnLWch
xhBIIBIabyTxKOw0Um/RrfdkqpGYztggBCR8buDBrtfNNMpz8ucAVsdb70if99JW8omkVEMbUbSP
l4kf7PEevGbC+Z3GEHpREST/DPjfSDG/H25j16CuSbuPSOFYitNggSKB3mCYDoR0+47S5hIWD7Zk
vrImT7cELOVnLF8NqzU6izkRCImaEEmNGakrP5WzkZ8whfAJc+JUKj58cgNXtnvvPPZ/pYgldqqQ
AOo3C69dQApTUFnFo5pSs6vJROIFYYvHw2xGWG9aTjh8K7uF969u68V/W408YFnehgquoKK2hFj/
1I9nTdE6hvhGH9vsBMqgeDMn79jvU6s11C8ZeJWffo3sdFwhJ5D0y2kzBRo2u+Eh69D+ImrJTMgx
ETgl59JBHEqxaImP9cbI4hoHfRGKYVVU1q6ht+UEpoP2V8NpRoO2IbdYu5S9Ov/T+VerYeLP1ttJ
xcLdC53/AizYx4px1Jvr7L15Kl9dRQaP7ERrgH3uX/hsycXlXitwfy8Vz+ETab2hNZXDhzXhpTBl
0PdJv54kN6KvmVLl6VhqhqzI4XuhrctnQpteTpa6osRSGP1OaBZI5bZusxnCejpA2Onpq6hI5in/
3/V/i+nWwm6NpXs1hCLq8xlOvsBnTi3UDhe7RWqul/VzChAZnXTSK1E7bQfVs/oiuF4ei5Y0DdM4
OQmBBBWd1VVR/IxtRwJWu00V5TOKuf/VNwbZOUudx3T6WMi5KCUTX94lcrUJA57b18wqIXKSV3zQ
JGI86NG4MFSmKCngmHhgoKuLHzlwEqZKKSXdeW6OalzxSErPKQjUKVZRVwwqIIE8yD8ANufwhvrs
komIV4BLUdQSTnKDEAtSPO7qS3RxGoVS8cQEFg6dFlf3m2jHvDRjpGKYsJLvBEouUUUUAtIc9ohZ
kY5A6mDJkI0C75S9Ie0+/f1dIB5ByNBzywYTIx8dxTZ+qGVkHuAdCuFB1HHgIEFDzrZl2hL3ekUR
jZOoOLyQuTYcFsod5uuV2eGxrl5UmpqO31bsFfh4R0b6uD8Axs7pp3D81JzZvJwNPJMcJzpYGL3h
Ci1mBMPZn1lkP7GfqFF+iNipawe2Y6xRajrrt6Vv1gSHUxnycdcx1VUY+gn+ntv9iWaXHLFckHKZ
nQIXAQWTBmn4fniILjjgjWvowY5IQFaBja4dJVC3UC8wQA2PqkA/m16l/Jfzndy89IXpoJ35dHd5
Z7Sm2bRtDNM4DWtiGHPJcb4cvkoz5b1+3kbRKoMOm7zPHJIAXxe7AvZrn7yYsohTdpHl5PyykrV9
rS4YoIUDxjC/QFRA+9qvmT+PEGzrvrLkw7cvqcpLB8S4pvX54k9gIelzk+3wLrDmTuvDqcbXUw6k
cIujS5SBwniJZA3aF366t2HYolszvjkTXYukLgoQhVdRCs8bfcTa4X0KwYeyGnLzyAZ+m9lGhaso
Mvt21AZewOUdwtnHzurGqVqYRa/Pzm7w+khWzosAy5P/EMtiaDF16KyreDv86MgaVTTxdcPlhW4L
/nTqnPBPCbvAZ9S/Olgnah3uoRVBZG/7onxxbXSIdP9cr9t4wAc5TfeDZvpuPo1Xh4lBDB7eoc3h
igoPwZM+801a3ZfurNh/YCieih/7xUWv96A7Xip8pICaumwRWw1x/EwX09ipeo3sxkTXBRZZYopL
rLNMZtT/lzCj/IV3GLy7DBTLz7wGW933xLoMddYxFpOIDZXTCOh+vxIZR1tw6kvGjHU/db+X1X8a
Gpc4MWsEQr49l+ktU7YQwmSrvkyPa9w2XSlk+yOxyAh3+YvbSqQ9A6phyjRjZbi0VxYOmHQe3w78
ZDKwLABBEGo+Zfc8tZkDtId3Kf3pj66o7qL/ttpLsu71BeSfs64XmSKFSlDvwnUeuE/JJ6Xone3V
VJVud523a3FCuRFfT9aMO82Nv0iqC9cXwisOq5ZXiTGZJJnujD+NunegMFVJtDVWHtpGAMzWPvJC
+5vwtcGcTCb7tP/SfCRd4g7cLfbQxtEPdFx83pj0lcm5LVqubDFWnUjKNBazqNd29/rFxi5tymja
8cjRLo71T7fsyvXOa01xGrcN+2/qAqivDYyxhFqYR31guPK6qciKmPBcL2DGaQJhtfyZkCZeRA4h
5sf3fwi6cVsvEqfvbTbnNd7oyXtyiDneqmqRlsdsavRDNAmUzyrirRCZCSYF73WD78seH6kSkVTw
3ZbeyK+Jr/nobJlp+fNcyN9OH7J0NepDrt8BL5MZbfMt84Rp8XKhuw1u7D/SHfnRy0OFdilmmsE6
uKANvmERzh/jbOe2l2ZIHY3jtejhJQYMQdH+mhzWttMQ+7TidIINo/sVSgzSbayYVVnGxahR6svc
/eObiQSjDC5R0xg3UdGGYNaBC+BIYszMZthIdGDAxZ0ZkBhA7dlO9+1+JRMa2HNUUzp1OedKqFgz
o6PVkUnBkn9cLDPZHMiR67N3OqOdEMMMIWfcgMpeX75S06ImFYQ4O3OzyC3YnVEMj7ej/b1eMGJE
9UN/TbXfUYmtIVUC/J4yFvX4ngsLCB8ixGnVMT3AHV2zQNj0UyCN77BRca3++KKmIrdMZsAJLxrh
L3yjk1aZlIJ4Cx0JMxWZGrcNiehQJR64b+fdTN+UCgbFJngA0NUsgECfr7oqKAaFLi9bYFpKziKY
sIes1zQQTwkW9vDjtAuvwUnvs57IKw/gUT+pdNBfXYaxMXgiU7moJ/XHpGvm7NF/jaSMmq6grW+A
ESBhO2bSFkoD+4Bp75m+K4ENt9jh9h+FOVNSLza6yCU/2E/w2qGXhtOtcKrWYo2tSn/lgzLQJij1
C03Tmq7WuwMudIS/A+wXtW7YAww6UpoDee6xu4MBIp6E3yr3U8dv6YbK8N/z8dQaVR82q7Q9vmrr
KsGyT18wnmwqW1yabLzt4XhnSXUKPcCNSGyANnDMZmNOW2gRAUP37yrbrgJ/WHXL8xmudjQo2/hI
hsNUByqFeCtXifDLYRrlUcCEy+AtlFPxshvcBlKggY1D2rpk/KfkEtr58RmNQc6o+O2J2QvHFfRq
Gf+8j1Ca80pQcE/qPtmZzgs9nhqSMg9V2EJpQFigeXDkOzUAPxxBWPY8cRDDAmA1zp6PDtBn4Tih
0Z775Ph67YidqZUqnlrzQilm4XysKKQQTyJvnqnnghHdrekMawOES4PwjSkb0V8r2Cue0Q1jaJ7V
BJT9OidouCyvs7b65geTO8YvKleKMnEu70MQy3IiuT5SMLqYhj2WnDTqy/0p+SsihvM1BWmmlkeH
NcEq8uQBATCwTCUEtBMMvt/ATf72uUTtRaskpzis/aqYjjfkA1EeCCq+heiBFSFeIYdNvLtMHUN0
rk+oQTxD5Qx5FLrQsHojkpmPgBctxrXw6vtrEspptVQGz0yx0bqyj2omvTner0Mb6O+iyX+WDYfX
M0k2U/LdGGHVcAtCZ2ooenX0wTnpxveON5mKF24+jJC/9HIUH4PSjPEzeQ2ozprKN3ly8W4DQr3F
vb805pjXkMYdbvmRJF0Hyg21TE9XeqHlLAjlei6DXGyzUtMTcPx3jRLdKNZ1qOvrqqQ5zXizOoqr
wSa5vZiyG3DgwNK4ACjSnC95e3LZ8NEqYsVhUKkXZMT09NcGoso7jweneQegtA8XWt0zTB/WBVpW
u6iWRdOz3MoCAHoZAERgJYzL6uHU3gW2j3uI3uPrcnhX0su44Y5kNI0brF1XzsrNq8Mvjra96Guu
7d6PNGaBIVtS449+it2O0HHuDWnhPcBJfpvuwLRCXQ4mzgtLNVgZquRT9Utp6TJJ7sB3gldTJ89q
uBilENSrkl1T3MDbtL5oFYJlfdqZqeYjeojL2o0wZ5U78rquebfhRhNHvwmt7V7xOmHoEKPZzmKh
XPl/gNQSnXnaRqkG+4y6chhvGpoeMdJG4O0P4S/4QYSI5FUBEKGp0bP8jlCe2svF/S7LXPGSxHM+
OtNWDb3OEF2yPTnGFxvLEOvzATy2LqkKB/ZGhCoKvreBKeLwVg6ZQ/a2VMRabK9VDToHO1tr69jF
5RdcZs8U0AIJDhxyoOlpGfhHDN0+w6tqvHhCMtmexXfUAZiVChZVgpn8/VWexS17A4DA7zUT0h8b
V+wDmC3Z2HUC4umUSWB9TjRAqF9cZVKuAAeI3VQsPsCjdeobTMU+c+WNTBmSB9qT+4+7lEepp8RY
MEUpKdMi1i4pCMqgQs+Ai2Kxzqzqb5c0QH3GHiQ6ZhhLofeFClumxB4ovx24GOiACzfRHFnuX7G/
MvVOXm5C/sijDPbsZWMscmkEQSdx0AI+MCF/rAdoJJh6EacCloxI9npqeWcQYJuJ9ypU4FI7ij0I
VrtUgVjYsyD58kwbSMnq880Qz0eNnQJjLziSAB2/0057t+OQvx8s4fzY4JNCrDhxzd9lpiGIpHiv
0IXewKFs6BiZiyAmkeEPjPBfrL3G36Jo6INtFz+9TGYlQP1v9f4ZA/dCHh/fjmY4D2bWbQBatd3f
emmAirF7VDvGYb0Ug/+R+NswJitHk4kSL14AbfnqeM89jY9a3mnmB2a/22DgiBpH5OaTeW6YElbR
VLxewLbVCjlw/bQ/7VzNTgZnQLqOl7dcLfi85ofSLr6FzsiZEYANbEjzEEquINbxwchY/Nyoh/uO
+pOYsm2dKvJthyyBlOVO+sFpDCOoyy5FC1xp/urdkP16G1LQKDhB0njQcXLuDnRJt8/9OpRgI1GB
cvkW6FdrteZalgXhJZ1OIGc4iUqGcHB963H3wW3d5uujrnsegWzznYCovwJ65y1Tjg6ZoPyIvKco
biBHZGl2FKKrDT7SzATVqFSqpsZHOynDMG9yuqFExEAFUY+LYnCKiQPdV8yvBNMEdCpsDakGXmGF
WJTtier5nhgtCCko4bghIZVxj3x9LlkBthhsbhDr+EuVRsPBUpkPmttQqb0oMh9MzYHfj0oe+TXw
KGSp4vtUc5cut/9HvkO8wADm+L8OiQWxOlFcd+zliniXljvRUxRpGxLlBleVkchMkgI8rZKPZ5UW
u4rYAKTv2s7xgNbA9o4sNjQdQhGqlz5fcOURDOYgpPSyE52+BEIvPOgA6HK1qMh3Ed8WM3oExKTC
0IIObYntyOOMnCZxZgB9T9EuxpEBqoN8PhwsAPgY3UbY8MaJn1jgaduuJ6YJN3E9rctRweUbs5Es
TpvHMV81C5urI1ryy/Mk3mfvyycr+okiL6htQfizQxNRK+njMXLmpeiPhLgG40IqCxeePH70E6Eu
dNNNvfK0F3Wr9z0ljlfBOGly9mHi6B9Tw1Db1T/Dj8EYfbC0yZbHTbHeZ4TtzMecJChN/JK5kqh8
GAxvEkLcD3SZ31PBsxHZ+P0RijpLUarywB1yckd8gpeHgzL70rzLqU2Tintzp6w/hy6qCDYwpUIN
ADOX/5NUlD25HFVd4RDpPr4H9baxD7ahdgPd+FyJ5KEL9sB89VA03GFVQLplCTR8iAtz2WYK7/34
kL2jNQ0SBrGYp6SKvjt+eY/j3fmwktK3qGjJtUmNlQ+VInDIex8p74qaJLkbDrJnokIcFUI2l0Rm
1MI0OzDW2eOWhtk9a3zShEIu9zyCSPcwzAbCuss1CTsrkPwwZgJnpDTF2J2QTYb27fpo2696WMRB
HQq18++W6KhMt4v0r72L6ogjbsnPnh/E+rxjGOGL/w7egRpl8y5X/wVkwGAE4DPFNaPW+udCa+0g
hZzfu0nui/nNM8APa+1MzHGxAa1wGfEW/jWRsJriYq0l6zou3zG+ksd2at7nO4+g8SKnGQl+BW7+
oO0CiMQIDVAnuuTmJQQbhto9tY05qmDGUVB+ezC5c86/vN2UWOPeHDHZ7fGz4i9F9Qn3Akc7FgTA
6IJ2glQ7cvq0zhG2uUd3Sf4Gil8W7ygoRHnxYe1Gth7hR2kYInqLAhqqcB0ntVjk9et0kBbPu0Jl
GmIhrRPMezZFDDCgmGRpOSanO4SHWw/9k351locVSq8X207BSo0JOeFRz3GMGga/SpupNrYHoUQA
UmuBliS8KqLeBL8Ia9/1gqYektwgn6P5sIHg6skoeOZAJgofyzaHKgF3rOKcBpPfI+0O40ehqaHh
+Rlmkq+ZkDODV9LE7ExhgS0rC5Wy/io9aJUjq5nO0TBOmPfjPN8a5pDG+ogBHom1IGK6JoHSYrBX
wc4KdXwJqQDo7nbZM59ukYqntRIIfmPXfqNfJYjhcKYCyIDC5IIvtdyPEQfBFgupt5+eNSAPI84X
CqURWMD3cBPAQBrull3XD90GpIN7yEMTGTgqgStGLbQILPeHk7MBy4yEF67+GbnMw+/KO2m8wBCp
ibKDGzXkFIQtkvU/tbBmBD4tMfCFn0CTgkNc4ScFazk4VnkMPqB5o41QxgD841bG5BfNxtpDrzgF
SvofaqWo297lkH1HMes4RQACtygzOYAUqjRIFNgh+U6q+Fu4V4wcxY4FdFxe5v8zYyVrsA7YgKol
6UFifH76BSOAE8oaLCh9sZDI0khhyFZdwzYJzFwSocCdL+gxujp+JczBRNxwlCaPoBgcrx18MALT
gpgUpl8fkn7lgGqhp/rtBMO5ZATvxrwKqgRTf/MvVyw3Iqc3aEJ6kRCG0yrZEdhrAgnxHk9qv92p
4GM0pW7qAzyPEW4zHdVa4JDS9uCIQrR+fNwv8KSFIMtN9p0lUnz5VriPK1gG7IkxSTFrOjBu0VY2
sNghRKmwBjcpC3Asut5+WPtMSkuQd8rl4DcZH9cfHhznZGhTzDpHhnMxXYeDHElX0ByMQzxl7bvv
NMC/gHQc8YQYFiU8nUrLTo2ojH71x3p2OnMrJ3Mu4ZzqztnnDHzsVwqGrRag4Xj4Y78ho9X/aBE7
RghNgZHMxmgCNBXysNQ9L5PusnR908QTHKjIcg7qtFufAGMBayDJxwXeM43kWx7dQjOJFqNz5wGf
bqrCRemy1l/QTQGj405SdeqSmTb8FrmBwuDcH/qw5S2Cixe5VnOrZ6IOScYwBEpuXSnJRkP5HTwk
8B8jbp9GjB+WgJJwWWkcuhukLwp6mtjk2bxBuJGbaGNANHc/98s110qhkrjezniiALfHFh3cMXrc
RTzTmEydmeORpOw4u6GDMGpBtrcqEeBlbOM2CdMEppKRG9rxglJMHwgKWpeZoQduDZFO4r5wzRKZ
k+ZLc2w7rIYYe3I9mlqqBCLiNJsm/1Pj5L51i1eCQV8BZ+cRgWNRLxJtHoqwfM0ZcMY8u2ABQBsh
7Npq4Fij1pUa1UUl3GivJeWBLa7lpltE9uPSVR7y5+R2lXKKMP/7S3d+uCUYg4xnHRgLsaoJ7UTM
qYJQmzuLVSspUcvbL/751TSGtX/S20EGky4ARWfp0nAf6H8cpWdANcmkO8dGPiii4yQF6CyzJEHQ
mV8FARrUaxcvs6BnBohQFLBpfHyA/UP/C9KZ7c368/h1azXC1TDkrVxRxHKSijbhkIKY1kaP2lJO
4jDRzHNJB+7lfttEIxOIgiCqN+C+CZOaj5oq7L3FOSPMuDLLHooyoTsLUU3l2if2HV0ROQuJYKIH
7JPs8KPMjBhEg2eA3XqsKVdofptQN8VtTg7Nrkl5H+TS9w9F1TqTfq3gvYizvXA89zYif4sSakfR
6IHXYQGx1znJN0h054eF0QnTjZAAodFD/9x74UXAnvzrJVcRfP4oMCWZcL16GOQ0ROamdd0rDPv0
/HPQt/0jm4zXLGY2zvhE2uyD4gcWvHM+FH5kQ/ugSlcaiZU0CwnNv3FdegmgIIuOgjWXTByksbeA
rtvWzCupTiKupm/5hZDDTDcL6khgMFza9bhuv8AzaHK9rYtdPiPGN5IKV05Brw+hT20Sbpb+8M5z
DP1hIay4gADJtMJiDEkYQY4u+KmMOx0fmNMsIKyArn9FE4VoHkq+d7gTpYSwWeW1F3HbAZbayfTy
iE3q93iXEAaOa/tEP7Ai7b3jmjH/YkPjAkNzBLHx6aEDrxg67QfdqEI0h+wBKtT9EMsTE8VmrT03
VGovXkiWErD1MlqVvKCjO60A2teYH88vJjE8eeUgBkWxkukWdGWpzFi7O/x9nzb4/8EyJdglD+X+
6+p65XsDvHqYw1kRJPAdX3n9IcJWgCK+VIYY6d/DYWY3wdw3lDFxd5sPAYFL9ZmaCFQ0wrDBbsjO
/4cZeRtaekLqtR2K78yUJyXQrDuqypf6m5Mocuio8QBlY/HYu0vAC0q+POKGKTuPNpOVQdqhFFYl
0BCqY7NH6PbrRq6/ILURq62LKBW6z4BwRcir6zAH0bJBQjkT0DC9OZ9k/maVsjaYGcs855mKScTm
2b2ZARYp8U5i/L1tu7jAVhtGe5v+VTR+FGpCgQyOdqFbmeLw9OSjN/icmIsj3fqQ6XC+6DkVlsqP
jqpCcGPo9tOhi7o67ubJrzDEgPKlIXjLBHelUxQhA8QYM4gxdZHvN/YqvYnk5NS38H5jgAsfp2g/
QOfMnW2sUjxbIGh5Mr6Y4AFADZ3niyDViucRa3bE0QavheC5QIM9VNED7iiaHBfCPk8UQJlJ75Y4
tLP3pmT+uN2xU8S9P298gxHZ0wRbgJ7RdyvEuFptWc4W90osr0TTuGakvz2w1/T3j2SiJ2tlSsyQ
NqmcQiiJ8WaxS7SWKFsn3oyVXpmu7vlepgtv1WgMxsMmSLZEx1y1LhFBRXLebkq1oxBhL+leEcVU
nzYDwmD/il7dvvg5a6G7l6ScKzZvf8Nv+dmFOb4+YttrFbNxkRXIdmIe0pEWw4hOb5SemH2Zrkru
yLfBCquVS2bgQF7msMCvm+/4vdFKs5+0EVVRMBEAwKPcwuKBm0VYMxgTdKFXJq+n9j7G4+XbUEl0
qk4ASpKQyUFUebjUiiZXOUu32pukWLhnwUwg1fMre3iZ5ZyTU1M9I6Y23yqnloAtRtkhHrVYyjqY
d4QUQjdf+uDppXKI5eQfkv/FfkN1oc4whTppd9f2ufP3A0aTF5LmHx9/sazHgbP3IjfVqHzBFwi0
OS+zhsv4EE3Nj9yyacjJvVnzyUfRgEtW842zB0d29MyWaPtF0f6TyGYmkgq1SzW5bawlAv6riiUX
DgrwMe/LE0hQIRJMF6msfLrIyr9yzosjU0iE2oI0RspyTFaISitGMkW0vcRIgEMSsUINXl534QLs
eUGhJH8EoXRAnKidQarD94b7xu2qbJDrvIWnqq+JILlQCRIBM31qPoGxQbP12CwqbsE0SoZ/TpCo
U3rOromUxxkhXOQSKqjtN+ukyOxU+gfEhbV+vAKxEpupdrfDowd1L2KDlo9QqlPAXsktUrzwDVH7
XHMD4bafVZGO8oh9BlTwWFFztwLBA36G26mrCzpU6l1wxw60hvljGjYTiztmNaM0kuN9huxtLMzq
DLQKEHgWfNaJkTkAXFukrTkPDkTEH9l+kDLiNvreEV9hiUFYVvyR5T7LH/iEURsrsAmMCiGwCsoj
BEdI18VMlY6Dw3zt/iQFdQ4ZIaldgxlubMzAbQUNJtOiNrIPysVtpw/M2Megtf6/nYpMJOaHXpb5
RqinqpD7XBZhaZWk+pUz6RlfUaGe1ho//HGUzbR5eqCDfffT9gVF30izyH5lczIogUjKWPOoQJ0g
7+5Q9HR4X5q1cVyosTjde+wQvcENLh7dXshukgex45Q9/myOm2Svn4uZwpDNgxNov+xoFIDLCxa3
E1ndMaz1HsAjvcvP5vrbZTCGXGlB3lCDLkqxLHT6wzriQnFzECrI0pAbhMY9BJdohenPwkigSE9Z
BrtKxawsIKwvNiTJLuB0A4hnggJgqBZvkaTnnpX6niwHd8nAZEI44rOSA8DFsjJ4lHspQn1kcxKH
px5KpuRtVykBFhTECaVnpoICX+bhEfwIp6iPCvNmDLigzbpRWYfmQqtTE+bDZGMB6aL4qVc3Kgql
9IIh1zRHEzHnrjJP3eKkirBNOTnh4tu5a1pVbb7Qez3HYimNe587kXh2VMplAOyyW22ke8+jTzla
rJrBMwtiaP8uoPsD5yhZtdYR6nUQjiIbx4LTXaP1x5+mDFdZ00CDueEWNjrPTQQtdhsOvO1Qp7kI
hkesZZi1oALPzzfc7QI4db/qA9QJo4D8iJ3sQkUnK+eqXC33ZdyQot+oXeiyS0RWsLxiWmRXHpw3
cm81+/gqYEqDJlyAoDAS7D5FH5n6fihB2nLC0ZRcx0NJknoMbgrvqQy0RlkwicRg6uezwOWGr0NY
rvCv69C/kaFb4f/Dnn4dgRExhOCZLZcF//kX0EFSg6132VRtxFvKCERRkfxgXl58q7LbC5cMPhuj
a5MnAolC0i1rpyQR8g8eaVcFknxNWXXrtRGJerT4VyDT31DcrHurzO805LtTmaIpGx7fYeTs3Hnq
zk0Ps9aDfVWITR+m8YCRJK3/jkGBB2QsQUyKcIMMpTfUYt9RdvWrAI/te9S4Z6L3XFG3wE4cSzSU
+vONddiMgcI41Se6a4ZtlnZym4Fwwaw3ZhMOWfhYpv0xu+yENyBzYHj9joB6PyevjpYhU1NinNce
fdNDE6Npb4BAkHtNVtuCmc5T59KXblqWVPN472v0CqB5bz9QBw7eFWLBa8GGimiUKr7oi52ZLdhR
wKZnWA/K0F8RGP3O0xDx7iUviQl4n89b4R1VL2T/pJT4xR6i1Ake9w18HYO29QNu+rq5RP7N1o+g
envNqcl2ENZv2LHZqyxXDYLtRlkMD9X8X4RaPeiW/Ls01/9F9vxQqrpPnfZ8sVpO3YSK44Q38F5T
njlTN0PYJDDkMUFLqwKD0X93FXlbsHJ5fqVMXPzCBzgqbTsHEV+TV0C8f3hfsAlAltD7lIHLcwmo
tpJZpLUVZacJZuxKRREWv5KXoBSCNw9knaC9QpTfZ4x9cccQ0mEUnf9IkqviIuHm6PHOQ7boactA
5bnCb3qJOgsY37v1NeM/QN5plF7brEBJin4y5Qh2JJsSPIPQtKwVM9nid9HDV+e8HWyW2FJ+jmps
QZF+foSW63ylFrtlgUIs/xT9DDu/B8eYUFhTp8DXqOGytB0vdc0n6lYfpr7Q1n3D9lq94rxm9Gvo
w2rV6ifeHgaPMgGc5G4z42Boww2D1fsD2rEDt22UONVQxzHwNo/VhedPofOkBTtAcYMPVSvDDUEL
OoFmJskKJo+9yxV7fXC5SYotrK7XfO1/rQnsqZ7K0fRCUTyEaDBEYwRiLkM6B4HdzWuQMpT9lFJv
Eoyv0tVM5VLFH+NzMFFeQOsLkFxLNN2OvnJomX+d3xhZDM6E1G3iNHyI3j5eilMGWGQ+oRzl4O9e
0yPf86lO5e/t8C+R5Swa6144MCv0fCDumrrwEj+r9qaBy8mAmAjcxKx8rkTJkGQUVMqdgEb0rgQO
6HCIEwzIoBzypUcSbMyjlOLNzyOXux5AKGJTl5T2j0v25kYnlCr+6fHM7tSr9uP0uiLl5uuF+C7k
Iw9cRL/ujpljXDHwKp1bdXo5eApDGPnB0UuwxSwzXf2JVCGNe1CzBL4oedrpH/FzLgqZ+0WGg7+e
00KlENM6vSdXEBNJZorhtVvGF1ock/dOf5BevwFLejBX+J7VCzUZuMbwcCs78FWTbXAkiebUZOi8
8iyw2GFwza+mk9rtUBN077eOC1dRdeRJo+ICEptkeTDjfAd0pjnuUbd3LhnNIwWqR9/cW9opPBBh
HY2D1f+BIJRKPpNZeZ/4tT96gjmJ4afheuk2kIdLxKMxtpn9OroAEI3P/fZ59MdPv0fyiu4dmGKW
cFkTShNRXJQ1aUV6MFhpa5BjD8dvihr0eLDGHASjkpUVaC9KhK2wH/XSxwXBb/ouERWur58ZeI6J
H7WnDKun7Q2TdLs7VCgmls+MUeT16M4MosSVtjbNgEg7XxcuwEDOiZaLVeCpDIOP75bhiefZp6yH
bQA8g7Bn/s0kUe5sP2rkfyWAba2Yv9vC+fiu0dOh+RObfEx9H7mXHnxVEASveB0puVdJKfPg5vdh
7M+NhUTGlrPxUKT9yv0+DmfNXUMXWb0mzs1ZNSAzYKgcfsAo8ahaEjTcHE5ysWX+mut9JWD662+l
efiTd4V4DKBbrLJ4Yn3lRXF3liNNxJIj231wDgXou+0vjKrEjw0QF2uVlxoobrbwTyOLe6WXe3Xb
xeAUcq8yXIhX6IqAdFVLvcnJhFJwTs8gyGLI90mLMLZitOUILCGI/Hp1r/fgE5KXAzw2Ik6oGCwn
OVhmFcSctCQHp6r6Untt11HKHGvLVZW2viSW/U+pulLZSp2W6RKni9k6x5kKkJnxjUgM93zDchw6
YUHXnDyAF7/yRgzC+e/iVqNeqHxvIY137P6n2tOfvuDwJHt6CGL5a+ujMaSvsT0r4ZTM7qsbEImj
/4Qz2ELbYIrBygN6PvPvHJYd65XRXd5Zbft0pgzDEAUwH76u9+IPLaMdmi2WOU6slcLCjj+lAQtD
6uOa5+Aygg2ChQueY5mWQcdwCOUkgPSdfSG6hitgG7hwoZUlcI0ZP7g0orO8Jm4BEDegrv3m+YdJ
MWp1LkuceNeyWRm9dmULL1iHa93UfgAgM/utkLZvlnF1kPl0MsK4zXovtgT41POC3y50H1fDqb72
eVq2vHpdOhv9vQ567PKmp4Ym6jUJpgfeky1I9kZ8Z+jLF9bcfpglafyiYl1VG2wT94IVt0oR5LmD
ZpL0bAUUreJsWG/dY7tesmuKX83uUzZRQn45KLR7cp3mVQ+MOW38jQyCJvsfiPkhqB6wTfFG306E
ppuKyfcX3TXZwCDGZC5CbbirnWhZ/x9oc7M3X3WvuNK4WXXJPzRdHFlJQ6d+rN0RUYrclTKXlkHi
ETO4u0pdgmnEWkL5w/yT0pwIuZ7HFCLrSqwZN8umd3vQMvz3QeLUR5SUQy6iOpHbLruPkWKS+hre
1R99xLyzYet+uFphjPbX7P4M23UhuXh58mbmnQV7SPWiFVLNkAA33C5axZW8jSkaLk0Pm32n7zP2
m15zh28ZNAfp7Owrvhwc3SkAEXw8VbqWfzGtOvie1rOIeanHwRVYYtDtEM+D1qeT0Nmq/wpasQQi
yuX0y+qks6dcxCi7kygUmMAJwY9XIVl9hmx1kRvWyyu9Nus7l3pzz6qeEQO7vCZhVDfmVbaXFh3H
qaXRSqLPcBR3YhiIZ5gaqqUD2o7ywEDGEW2ipzM6wfeKCnWdNc5lpEtMvWuv9/TqovvGHqCSgo0h
JxMH092dlDVa1KZ29tlj2y5ksSiMuAD1OE1xpUWhEPmML8Iz7Rhy+liify1VaxS0q8bA9nBgDXVD
U9XBirQb5+E6hrXpq5KH95fJrc36HEyIJaRixDTDDlfVeFPpUQ5wh9pNKDH3/Ullj3yk4CVrjM74
op60+CsilUjOFIIQaxCQRuBVNYhaZczl83+Eod4QxNaCl26HSbgfQ9CjOseW5POqjlvXaov30tXo
3sTCe2fYblngujUrlmmVriV1rS+gXzMaXBnT9KjtakJ3Tc0nrLtkN1IbM2gJ6EQApc2ZheJO54EI
sesnK72Ehg7JHVIQVP3hgVGHjygQUpda98dBkkSwvl6BUTF/cB5wYs6TRl8laEcYQUCrNH0SaGb6
+YJZKYLGpuf6V/PwewkPD71uIZZlpqKoQmFdbAiIkaYNgy94+6JAm+2kcTlkdN80xQHWNTy3+0Wz
WIdmuXk+670IH6ozaO+fJzsJ5/UOrR6yRwjMzlFzMqyz9mjUOnbYykPyd1IdKhnpJ4p9wOaAm040
lEVX+Nj/Oo1+vLR/SCs934ylm+/NVyGgnKGg450rOVqHtUEkW3DvqDfk0s8mdyLcJxzdL8ZWpA1k
kIbaQbSY8ebSNabyphuGkOyPwJF8aule3nOKkT53tqcvDHBn1X+vIEa6AdG+OiG/4JFu/Y9xYGnN
Fc1Fr8G6dToA31QTHtySQlkvByalhFq5+fn4hnitrXxg5jaeI5C/Ne71VeRwzlfnckjauBaVuuY8
uEc2aRB3yofsPr1ZHKRdI+F8ssJKHr5mJp0Q7tKoug00AWkpirVASRDDn9uvUi5plY042x1Pk7dF
rDKF0HKgOJDVw/VfEYzv5EmvomAA+XN7j4UAhojjWaZ1KeSBrCQ9UCVdkS6JoDmrNBhoMyxuluQf
RHUOOhXrvnfRIbl5Q4wF8S2FgpGB6bHXHYWX617waIDXyP0zjqCaI7E1MPn60Iinj788ZgjF58EM
C4Cg1jsSFlSumJPHytbtz0wva4Gd0KJp1tnov5W97nmq5KNwrzyAmwSdSBgNuNF3l1ImiL78Cqdj
Wr8ilm+AgMpNQI6S9RCs2nx1dUfN3D+dyv4lkgYdod6g8ZtGan2ItnJIzxVFwZowXM1mzIHpygH/
qjX3I6wfttcA0MJ7123bQJqJVgd8/UlSwCY2Ep0eXkiy18bhvAtDqVNe6vgw31uGJQPcL8I0LIHT
xWwR/sL2XFp0oAFt8la1V3gfOa4yLGev74B7UFann16xB3xWgv4HEHIdNWApfcBgHUOSCv3ud0sb
+kJjY+41kxliQ8vRRstvmcGh5fxD7jqIZGMssty+wK5B++OWDnXPv2kgSHS52jtbpnNGKNzaCFAx
No9mlp7FxPz8yCrK3IJSITn/euHL1u0G+GPLyIayZ+/mbuTgLDOVL5B/cJprHf5O7GsC+tWCqQ+S
I9K2e8sWA9lRXXrl94wM4WE0wX9LoWwuvD5JWoFp0YyT8sYKBZw3lGf6O5IwLoaA3D28m9Ys9oIF
L7lrtT3yrsRXy+VQVYA3K4mMCABFprOiEXTftz+3kZ63/y7k4GRIcZa6V+yYiUoY7vgZ/JoeuzDu
CR3b68CYR6RFWGY/TuOcRt8TyPOarI8V064yxj2qr/no9/PM/+HcnyrTSrWwJiWj1Ky6lrP8wfyc
vOL4DXtQFzNpJq19403YGNAWYbLxoTuEElkXenxOV5XxLB0EFvrtJHeya15Bn60bqCWdy9qUX6dM
Er9OT8GX6AE1UyW5BiIpnTewjaSneJCJ0wLO+QZ47pKU6m271LdFqsPgREQA1nYBsVxkeLssy0DQ
lSnBXXDTtAk2GedXDJRzkuZuVoES3mEYF6SDGALaBXDoCeYZcc4lYH2WwD7GgjIPKDvqbulE/e4a
wbO05F2DT/skInUNRwW7mHnsGLZ2TBwhcqhmNsUUseCiD4Rb/BkzaBMpIw0cw+Mbq9reSl38DUAh
SyeN1UlD2M5NF7wp2eBzeh1kl2rNFmIY1hwHRfrDxLGq80OWIWBMrncnKGmXc5yB/u+MaQ3sRX+s
RMonPmjT5ACJvZ2vRnkRm3a32g6dJzR4ZpZ1q3EyjF4mPdPxitKdUZt2HQ9Q1Srz7R0S0KHk+lxA
3OgyZH88FHCER7V3uZwh3o9yYKcXOjKOq/UVI8FBKNd7VcYM8Xfg4O2G2LuPRJyz2rtusf/haCGE
qS+gCRKgCfWyWr7vauswYLCoyQtUBU/l5SWJgWV6DPg0NGdk+ncN7f8zKTu3yLeTbc1zNRddWgXX
RpnphDJhlUyIotTvmHgC0D3Wr84D+HNQ+sU7k1pd1R8GCntMJT3fL3BJegSiQwhci8KPM4QTTkFE
T6sgnzwjN4h3xK3Stiuz2rOeMkH7DlOurUxGY4cxZPzNrQ2fzETKmiU/1kNFAJpUSA30WpOeGgNF
gjdY1j/5W4yzqW2WV8wUvm5KYc70OL7v4IlavMngBdUG9xh8rSoLtUggzGfgd+Bhcy766HEvZIdv
+7pmovhubSUOHZYy+vFERaQsyeYt+qU+klC+B0a1p1jv29WJ3UUsYyPU7UzsdKFuh+Hgf+gcakuO
FiDhePWDYdybI7Cex0b4U3d+wbdfOy6yUv0zQgfv8KY1H/vA9ij2dxk/ZicIGaxUwaBfX2l20XcA
Ek7l1WkKtMPlrmK92wibKOkJJ8DhkvsU7aGSzN0RSxReH7ugBzbG0nagrqjQ4v5a+BBZR3qR56zf
55VwZ5UAPtumE8KQCdQCe5rs65OIlnQe7cpXuHmXNmh3hC3HRY2cdXamdMOLHZHmZlkE4pVkYAnE
gYg67Jwhsp5gd2QU+CQEHZFAIXA8gYi5hyHNO1pUAbABctzdqhql5MdDicxZCh+4ybQLYt8Q/IAL
2yBQD9FrTUzxft05pt2binqLvh3pacY97pVdL1aEP+w27CEGs8gFWVDyVaz920xbxBCaaG0Cnr7S
61IlB4l7LYo7EY4m6C9S1uRbbv7m2kn9cVORAdZbrmLB7/0xHBEhwEX7syompOw2yhUkR9oR95ua
YJ4JYuxyfvPtSwjPZDW0vAJD5KGR59h2R0TeFYwI6Xg88vumKsvLSCTYIj2tKKhABW2FaxemZiY7
Cx/E7bJlRIS8VwUk3LEYLFNAUyI6N1BQenZQKYRn5G/uv/18thtJx+s6gzXtZiertDObbyd92N/4
j+0dn9HAVYIZZHnuxXb++vQxMXGeS7vR23tr+ZOzFQvBSH1aUwW62CmsfcBlGYzYlr6c/6wVcR5W
LmnIEtmhmVQDvFfgcCz5WSibJtpPI/Q01KAHYHoBCyMI6aNW6FZrGS4b5lIuSOR2Iqao6175C3jS
cdJuHzPwDOxOcH/0QK6KwROT0ZxsjZgHij9wZ/TAUkfUk7UoDvyUSlwV0zcdIQpd8j34meyIsqOW
n7mVEMCDc8fKpsj+08Zn1zOpAa9PhbnK3OtZ60qw1Gdl1F2b2Bo0t+cvPZAJ57C5V3ACgOnEM4Jw
J6nBawHuFJe+3btkfRwJCdMOF+RKqUL6/NsfijoZkfR0XytbQ9w29og54Vs+y3FtbhFHEluyaGQJ
gjs34w0vSp5qNTLUCpFZLXmLEapUK+kX8E9uqttUa3Mzg9Lwrn+bfyOYjkK0dyk2yrPehhbP6sNp
CyXX4t9bS/nePWPko66tV4QwCgcqoKCP8DEm9JNElp7VqtR9SHn6y68RsnKTGkGkXvll22EmG0nc
HWXrauHvfTEQ7ZHpZuhGrpd+3Viots3LmkgiGV2fQFUHOgxFqF4mnvsvycsO4xf9HcWqa26E6Z30
eI7Hckgs0ENClNFY4MwzqPYfefAZIVXkXlyapHdMaOts+7St3LbWa7xwSKW35dKZvJQgr5FHY0Ns
M0yt+XD5YqD3wFCjvMZPUhr87jI5Fl1pMVOuYQ22l8pt6SFrk0YRCl2hpg8ZWriCJxyaU7NUTu+j
CvhTJhVTxMloK1svrgcbvzF8brZVt4zwxOn6PEn8WWv9WY6qM54MRkkn/k7+UF2KtQWulmE4a82x
Cp72mTV1Ljwrktca0RB2w3+KB4MIlG11Q99JIETOC20nVnI3ozOlqHpttYhfOZZPvyeNXV4a2U3h
b6hb8eLW5YB7QgTAAOCoE5dQUWqvXrg0z7vGgZEJokGZx/ngnFp97+NmC1CvqBfhT9+G4qHQkFpM
1id10YQ30RH3WrVRKMCBlKm+aF27DpolvbQVKm5NBpWslSJZF3JqCiu22Ua9qe/IW/EDuErkPnIo
VgGkgjJ7KxI+V/vFaehjqg5NmQpqLiSC3rHJ6FuNBT6ahg+ZyaXCtNJ9WsB/Vxz9U6idGhr8jc31
DfhBB0ppH1s9xhFnE5cF5G8LZn7KMa1vxQ0uPkaOvOFX1P4RvddZa6YwLirRrbgeolrFMz/tue3Q
VOsGOFNcO6MQmXE7DkivzRLB7PjCdjHnbmE4QUmH2MGsBrS07ILNLKNA3nElJADoFGtG8anU5NbG
fQsL+vR/HGa/CaC8WfN7+JoPeCEOSibNd6L7/1UpjbXi8MUrcs+6sNHpFhKvuI876k4rjVFnaT9K
eL83mfQ/lqpU0u8Rys1zDev8hAVK9xD8VRY/kQOpkQaQ5mMKRI76euSw/8vXlW3C0wFyu05n6mW0
zGYMC9KJk7OHFJYr4F+hShGmmQqlkhyDngPupaukz5lqszD5+6S7qzjaOLmkrrUVAossTyY+HEU/
MWnSa96wLXuEl1gVC3ujUMvQtXDvSc8D24bI4kXpgGXOR9hW4V3dr4yQLEBLqg/59oUQrFBa1FsO
gibV4t4Hjnh0ymIAhHwuCpZ4setQYcNXFILzRGLTFJVpoacDzXHBy1/97r+zsr4Sihy8Ygvef9qm
c3vQJXUxv61sjxHUaPpJ9F6v5ufTUDaqvBuZcG2If5zFwLh02avKgECN83j1hIAD8xPW+Qv7MGIi
nom6tMolGheE7u9+1O3esxdEYkMWxgRwypdw/tvsO/WXn0GxQp6PI28Y66sgzVVz5oLMdz1sId97
UR2FZDOwIlDWIL0sYQg0EDE3e6eqgvk8AmRl0ch320C82jM5O/uMq9xN21zeRuak9Hk/gw/GqQLU
mGFvlRft++lnUb+BY/imtzT/1N1U4RGX9ZQzaQVtYpKEN7JFOucuum9CVWmYZqK+Jaf4eEanFiwl
Y8shYp5xVWC8S7XUE/0sdE6BOyjDu1fcDNR63oJeXR8XhyzzPIsVOJdTs+uTEYz1TMhi/OCh0auO
E5fUTmeXjbKZlzKZGz1d6e9uWyQa9KigA0Wu5+5gwdPeksPg2+3lFgOF0LLlh6TJyWchUi2lWkG7
7OGSQ0mpooqyfuNvH/jXqyqdMA34p7geQT7lCjmvMh1myv9Wti+kO88sZWN0sE16ALq81y2lXbQ0
ruA5nfaJ12KgFBua4GcK8Y1KMRnBiS/1nmy8odCiVx9Sf8SF6S6tax9VZF7rOJHl0UzJTWRwPElJ
7PQX9wGb2l/49jlaUaK0fehuocskOdbxH5yogocanaCrzwzs8lfJfvhcert6fXomQBJsA85lvOEO
cDYYzrLTXQuvq88pj75TheG60F6SN6cV6PVs69as2GbSsytc5KrPL6MawG6AsaanXW1ZiPqlEwOG
kMcGKm4oo5fOSkpmITIpqISVxDtFCfg599rjoKBxwu30L8sA/Ry0dbMFhLPziUYbeT/D2wxfTKGU
TpRpDoAEbkUSAB3OqDJa/G6NYCEUQRukRS2jktfNOitlDWn5uFn0Gi3cu5AExNzq+UoekHC4rUv8
Qcn1gQZIjkx9CMw3yOrOMCQdfVizIFlVEk6wzBfjO1T6tDmokJMnlggS+Nw7E5e9Rj2LtGby2/Zi
JGeDjOnisX7Nzgb0rV4SLfu7QLVh9sONRvDg//rXDQyAvZBGGDPh4CM9OS9JYeDJWvuylO9efW70
rqeR0ip0CVUNfvKyv+4EZiSilHtPbciXkziq8C7b71hTEPy+0XIEjINFvVnXeyFT13eNCHyqsZ8l
mLsTY3s/tZpPrzybY32hM8TxVmX77t7TC/JkjI7QkEX58ifC8xCuITRxBh/S2cVoxhavObWKzhE6
vW54L9TBgDzeMW63U+mj2cKsfGQR5qPRRLtTYHTQjgZyMPL/s0gG6QweRdJYVFJVIXhzf+js5jnZ
4wA+5pLffygU/+R7CDxyciAqaM8VH8yjY9WJN4DmCt/tkEwGncPUZu6gg5lx16VHGwTRYhsqHgyb
waDppzTwVuWQPTkAUUBrRIgMhYkFN6r+l47q2BkMDKN3nqo2qxGomjQ1zS4sPCVTqPDZKkucesWH
zAx/HIw887ciVUTvs9f5A630DSGpjgmVh1HesZQxP66cYKc36JVTfIKIMdmXEEdpSvUbcoWyq7JH
EOxZ6Av6nGpwFVANPJXm/JtNoA8GeT31FZ156YUKYrnRcBVF1PWHAAD6+h0BSM681i3XuNm5yQF3
RofLfPMDMPBRRf/5Xf/O/2nofLUgY2E9jRLZZJBEAtbKG1fUFco7TTRvJOkpcscqDqq1s8Mwgs27
9F2y/mGJTUNCNZfeVd2esA0XJC9f72oTJwrbf52bv23IyjfFJp/PacCWkLZ74IZsxaPfa+85WK5Z
TU2dYIKBEVLhMNAN8Zzar+JVZ3fetOgw5qKwaIVnaZNGoNOTgtv8o8GlncCEb4yqX3+ZeH6t0Ykh
fIJ8Jj2f8nCdqScXgk4PcBtATVUKVPNDbT/PC3sT0Yp1NByh5Mny3jjZz8RgNkDGWCNFgF94ViJC
WoXeBVUKXZbKvJ4ma2HPqeGVTyyCdVs6P1TwEeb8P5Jw78hiSMckxpBWWQUEu8mMLCz0BWmIitew
LqvMFIwlDY4Nv4nVCKyEreRMJphHlXQ4CCRPGDVEo7nrrydpc7ICLB3MtypH75jGDrNa4Uhavm+J
NrRQNjhwqyDNsWa1DL/8Ti2qxBo+W7C6k9EwnncIbwc5uFQJ16db9UhkOwCjLljzoFEJSPDX+bCT
ztv8M+UtVFdn+qItDCdJoHcCcxTan19JDzOp7Hwqt8ObFK+Fsvr0ZpInJPz8JqAqwiN0TTlljD6/
TDefXkhwqYdjbV6l1kR5n4gZpyrrOSKy/3U2MtwQj1IOx4T1CixObys08zPqbOhrq83w7S5m949L
0jBoqQ7kMN2j71JwVhl0UvzIYrC8l/VdvH87CC+IDxU3yT0BEGkgrrmVsT++FFF3r8zq3om71mOS
pvBtmMC26okX9+amD0GeAkf15E/yxPZQ/dn3c3n2299hWlAKgPqtp6KwqvksPqCYofcnQRLpevyI
kxfXDeYhNq5VLR1bFBVLKyWRuMEQ+OcwXFawNCL+cwS2R8WikPfmrIZdpWxPDFWLF+32jf0mnfKW
i3+2WnzdIDiXRJYxyvo2q2pqbaw0+k46OZdRQU9PABM6qrVlxfneY61sFhHYl/NjoEmG3J5hKmJU
e1jl34SHs2PEwMnEhntNF8E1TSFw2zf2K+DYh4fj/t37vvdTTixh/qXohFegQXK7bgbr35py//Np
ZJF0soYGUPbAKygtylu/m/dt3jOv/EBsj4mq/JZTZ+wZ0MT4kLZFOk+6BKXaFW85e5MF4qSr89Ya
6m2NsDfxPS9PJRcbughyjTQkygF+bhljoMpAF7hTCT5N/oS9wkEoxof8Z6r2Qoq3ZHvRVAAJuVZQ
zHlE9bGVtHw+HsGY1VSk5WltMA+Q2AfYE+HUnN2Jl6e3bQkNg7go0DIPSwVzMrSbgG8KocrO+zpD
r0c6/vow2++nFVL7dVEne69z7ZbyKiP1q97ayI/4Xj0iGN2m7UEOc30/7nP8T56Cprb6c0KIkt0B
dw9txglQZY8sektt4jEtv7rQ/5CMYHMPd6jq8ziAil0LfhRUCglq8Buc2OyiSuIz2qwpuvVGtSjX
0VbjKEAHztw5/jDlB3D0G/kLJU6hyWZ5jtEHZuPUSeLZEdTuX5UyjSs4pyug91C2xwddS1bWfyqa
6nG/s6Uz3IGBHt0cYHXv+txoH1jyBJ6KtMaxoYodfngjsMxuw+HrHm5UdPoYe6eSjEFayKxafeMU
5jMmrYgjgg4q44JTI8or9RJfWd2zydPHWpBA51aG1OyLRYDbNf4aeUZBEL8t6Qoym5Xu4Ingplxp
XBBh42CFMTcx01EMczz+AZOTTsAfRr5kAIY97eBsP1F+/q7AZnPZ5TR7WHQ5up3F1c7pzrMet9M/
OyPVrJYSk8xO77K8NHxTgHfWlxX4KUjGDSDLXrf/CBDM0eQGcvSMO6iT08n8EGpbCGlXAVz8JJwR
5MqbytN5MnLJGuUrI46tA/xA4p/OvBM8zbzFzR2pqA2J6pC1rDYcGr4i3lSWNG2gGpykbV1GVdHp
dCW7zvFjMBJuJz7+wyZiTp+zKKU9iIq+JYbQ+ZE1vvNh5llnDBCrvR0MqwU3xQZcR/Nr3KyFcHb6
TsBzgFdli/rn3kiXCMSUW443igNCDbLo0l7UNA5+vAs8SfXs+tz+BUYa+/Hq5FtUNNhz6jL2uH/6
TdCFvCDqbIcjrXwQRXCsTzFCybIulNDTbI1lWnirTpdEMk7lT+b3mFA2X5gn3GZsHuWfFcVTBKdx
bnfN9kejDvfk2u0/5hXf6dh2/0u1B/6ZbuF8XJyzBuuasUXThsJKKGCPXtlbEPAOUD+QJE0K+3Py
bCbzZNNkTw6YaB0h3qqFxthULjcBqDRVWiTbkRZ4u2x1vUJKMCIaGQa+EFT52RIr4r9yZtHECJ5q
JUcUZ6paApXHKHMNXzORNmSEdH9p+u2ckMW0OiGYjw7OHBPd86Zulr563TRs73A/Nf56XQokS1g3
FtOwW7IEE7Z/1ST551J+3jLqA/MdG27oTIFlB+fp+s1H5nj9wPJJPMvq1HtJKjG49y8ifj/gZZLu
Qs/2GxL8YkVZnIO4NAjyj7ZP/53Fvp50N7+zTJZRMY9zS6GoYiTASwkiRABM++QR3ZaRaMv75ttF
Y+he+QhWvePAENDJIMn7mPq/Q2MKmTIm8eFOj8nCSm7rZGXjgU1mSgFB8blxFf5+ea2THO8K8qF5
zufKqh/qYZbQ/t9+c5HuE5VRYGf0mAPvtpbTVNJouxu6GE7aWnT79jFiGyZAx4LXRsK5UoWJgULs
1RsryjQFRhfbWrYnYhv2OdGErIk72T97bcoZzhX+xluMcCxU1eYPyXZXADpfC6kNAOw5Bf6QW3Ka
J8QXY2zeYAh77Q0ULT45Hu1Xqk8n2SCVe1oy2fOTQqrOLOleU1tQPOmL/gAzXZNNRZMInIG0lBJt
RWRW45mf9zdtYWWbGYOD48i3yD+y1i6dfzzVdb0ESfLJtZo1ZJH+fmKuwa+jDTNmsMRzDAdFpOCW
Daa6JaQN9j6xKJqXsXzwHJ71KC9BarLLza23j26EaDxgQ0d/ydazzzw6iYWIzy4bJGu1W5QxdHDR
KIv+/Pi+30C51zlbjTFDEICg4PQydBbSPMiHm7+VwBjcKq9j5Fwp/TtX/rC86/HykZXP0+lxPp6V
NmGm8qxFqRJhttrlcACGJhNG8gFWP1ypEW3yHFkx7wafoXOesGmcEAR6w2FfznM0PGsqd/thnQTv
2EsbYf/ns9OjB3SrqFok6k64H7PMrC4BDNXdgZVwlbZU1uIIIUjIMu5UrwzSq5DgNHcljiWNbUQ5
NT5XxkUVRoAG34A8Sj3l8gtY6a+TIEi/oNW86YnjEIdCkL6DaWAPs6DSxkkLqLPxgV6KJw4MHXkF
q8ZB+2dRWpZ+fUmp5CHddh9l4sWceSd3uDYBNdLDT3MT/h3M23TlpCfmSJya1FCWHaKGf2XI1ehG
MkFU8IUQLLVbknoUTKzW6FdQkKshiKjebcu8rxVxJNdb4eFufiWWPvF1f3mUnbax/kYbqT4Xbhut
Mnb9kYUlKjR7etV0yubxZk1RP0inqUF+SJVFfOvlqcjAmUKWhRiA6caa3N95eVfOQu5EFWBdi/Tz
M4iHhorAzx2N9TdVGWMYqIQOSibrmrEucVo6UOXAIhfJxgSILKQ8lO6hnCWLmP2i3XGgcn6W0+f3
joDyfxWxXuiG/6mbKMEqF6B+QzaFCSnNTOnb8XqcdG6anU8iJ7FAcsHc9+JCSfmuQWLzQVInyAAk
KmoDdcUAJPljZzXjUX2RWLHRMHLbEhrEQfbfmJ+NbLNIp13qfR0vC2wsewczDlDJ852TpKa4HbyM
jz/s1ZT34N26JzqYXykLa/ZPDZfX5faUZaMzLYfT4fsHTcTXSA22osblyJFYP2gBiWrh9Bl/XQ+8
7UETFRywd8qSKVj+2oJMHMlQy9606KTZNGTbEtOKLjen26TW9JTiQyYhvWDCLzdqiDMeS5y1bJMs
AOOc4jTElro9CjtctY8JHzk/o30JS06CqwauTjLzDdY801vr+TNDKWRRwflQms8A54S3Chh2HF6A
xckTi8r3cFcOL9wyaT9TpZsGg2aIUx6CgWr6G2NEsbdYLlBTPJpRIjTHV/SuUyuwad2eCnhGflrc
Vy6QBjafeY/1nKksDR8UZYtCMlLWKxsHcBCHxphiUmJcCU3jQls0TMgNj3S7LHEGvw+vLSD754/G
ADOZT6wNWm/pKMBdtl/rp0UrP9SbMVMy85qNkwX8drCi1/3d7287f2vOqWpahiAw+xaW+vOyV/lf
+wtA5tMF25jJCtPJCtnCLzE0i3VRTbRGlGRkkAcvKQNjM9aPbyYbFa3E3RFNnnqszE2skMvt/1pg
wK7F6sSpepSYoM8tUqZL10u+nyS8rYAD1AcDO/X0nOd2u8QMrOk9hCn6g+hbcfg4RlnLpCKHmC77
B88023nJACwEdWdYExGxGzshK3lPf73WihrP/3sRg5aH7JhG+HGpZWzAsfOA5TIY1x7pJdLm5Adp
z3ZygxQ4C9RYQyFiAAmzPFlbUmgfs2ZygSE9mvxotyMI5MrhYT1dX7Br8UXmWZW24wWGpZbJGLwS
B40VVqoXUhhNe3vTigWvqzIcTw6t2dZ97pfaOD+IH1LdYnPI0fQEfs1T5wisetpRbuqK/ZUmgd+k
xHtR5cR0CM7Yx/m26yv0B+nnkfGqZrBnUGSGSnPprsMbLVmKiVVgPTDYn1P3m0amX9aLONUZJ6bD
XXyyMZROzRaewZ7Q/xQI67CENUiqRp/JHH4ZkzL12TYbsqjgZKcq6yPYw/+3twPj8ZcmSKCvVvhs
v6qX/IwjcO5HvGwphXZNZrvaFxm5+SUeiJZ+qJxfTH5lqFueftWMl3cqX0VpkVzeTSRXu40fOenn
lylbn3YJhQoNk+I99NI78Bwo+SDyZLhehEL2H474SKkgn6ghWhKAX8ehsTbfzSoNDDF2MpGtNs5c
n5o1/tshEk58veMcNQftmgl0BQaT8TcnHJ5NM/5PUwqzAX1QRjer1Ni4KjzQeXzvV35h/G28DCsD
zWgvi/PasZ0WSlnleTTmpOtwJVDDtO0tH9WIQKVmSHOVq8z2RrB/mkHXLuAtcIHR6b0FcuhfoAgt
lXZBiDgsiadHq+MBDZNhcIhS3cQy9eAI9UNk/GV5meHYdOX/BhHi6oVKpxSxsH17pB4nowCLQmtf
+KOLo07YMtOliUAMlai0Ug419oh8NWdyCRybcQo0FKGtXH6vxLj/HplnQQZj9FcCRjdAI/uYO1X1
i47UA6YyYjL9deiu/E2OsiXm19ec6eflMPYCH+323rXlrmiF7Ks2h2prcrENivsB4vDLAjYkZcLl
014GOJ5/Wu1Cgti/dkFA6exWnowVDJAeFXmMeE/8AcVp3S+HiXkiGFNkSWZADylhNAx72jjcFNxc
uwKSQaBVHl7+a58im0dvIwfi5QBvVI1Ro1SmGlSBbfGXjjGjBruUCQwsqJdqgxH50Lo/bRX9vnn9
8E0wo7FGEoxNbJoH8owBJ0DTigzkwT0fgn2UYFZWijJ/Z3uuNp2NYixFtLZGI/pZi8O/VOn9BKag
hel/oC0nFac/7YcnWT7w7AtdkC8DbUqc5MGDrnryVGZyQZtT2q9xMtDH7omOnJIWiOFnLwWs4Fxc
W6VmWeaR73yDHnLHSMpYD8IDIGOHpy89H3Yp8IYzi8t2blGx+nFl+S9nNHbDwAn2Yh+dilQaI20n
YzmAOf6b0S7k3rlMgm5CuPmQspar5tLwTBUQ1u2vrnLiVg/56TgkneioiOIdBpNl60FsLemFL2R3
7FbGBa1VJnZkjluHcEPy2FqIsudS1Jx9ZaN3T3pihqoyu8mWYExEWm47YpFKdf8k+zGUVTh65R2M
PvpF2DWRZsxZWc3MWObkLlf8rcDamW4FHia0bQQuv6o0AxRekFK6JITqNLElrHgJNQf5azyAy8Ad
erw9s6teqtlnKCXAe+crr6F4/Vuee470pmRegU3OxaS64Er24Mgsz+/k1ORoo5KClYAuoTfccr3P
e6mnxQqTfftNz/4edxyW3bz8JItMrfMorrU6GQ8ik5d20FYqDq5O568E7hCXpegnfRgd/iFr9rpl
935p+RaKG44NcbQ254M4GVismINUzsOlVxQvkvwjkEXLzxLr9MCoEgDleDUoujQ2GlqEG9qqWjdZ
8dkQjheWo9K9KWBx7h5Gv8H1TePrWdgGGtv9QRjV2BzwdgTe8XCQIYJiyg+6JRH2pMiQ8hs0Rbgu
5PflPN/EHb/cAI12NWNo74jkRCyOIWTw/Ns7yreZBQnCJPJzgdawtxsIa3IU9NeGkrqlT8S89h8r
javsHi4qvZ8nYuST4LwB8u4PY787QTuNnQXqHSoNms+yTHo279lNqKYtcvbpHqEv2OkvnhZldQlJ
rAfDsUnozhYPl6q1ex7rw1pzUvDM3+AsExLl3da3IjlCJOVG+LVROT+eFvypr8YTkZfLqB1h0XuZ
GKlvDUKBNeXZ+5GlRmugs3j/giJ6OdV0fZQ08TFUK33F8sOBNECb7BZhc0ZboLbn8dj2bHzbXaxy
K+ust5vs0vzyRDMa0YbuBWUV5+nuRxS0WjdI015qP8ka/EigY2qRDTJT+MrQAN/6rSeWfu1SgL3W
E4eiFXeI6L6kYwG87B1ebQDg7kpEZHdwAn5rNWoehkQ52vAdOMc1VuT/5Uz/JspDPC1+iOfYC2+7
gySSpk5OOmbj9cilC2k/lEmZ/fZWwsjhWKC41hBY3S3HAwCBvIBVl6jPpSCyR0jt0jcS2SJaLLE5
/fT1BDhHhRYkAoHyQhYpXH3MRM4nT7h7r4AuwAysqVSVkON8I2CMGtv0v6QS7rhjn/Gg+Ozb/3KO
DjiYXRhgdenRXK66TOHiAa8Dg6LvkxTh78Yq96JmUWmhRd6G0kSRwucQuH+RFLpYn5W8ACTbjKLl
OWj4QG/QeIpTg7hKkyZmLX1PwxCwoO10+7OQp5PnfCAmmFGYXTYM4gj26tfahKsqSfAyQHBSq4GM
W4BKesc/7laFJpTWtVFOOE4xs7eKvf4pKv3iiijQ61cMk3IbBrlKXSDZz2oeG3P8qXFZwy08vAR7
4qGlW8hhNKqEWSgJKBUVKjRKwdXXmzw2biPULnYCNoHS0HX1fi1JDEE+HaysCNXztZCBw1Ca5ufL
3ZvQkUSBm9/fSa++8fOo89qt2N1UosBqj/ofZpl1ktdkfM7sONeBGtHybgAyyGOmsl1Mhv2/wC8K
4rqAAXr9q+NRUKTcbIQSuUX/Ri0+Qvgs4yf1gwVynM9t5DFdtP75HmtFxuAuslRLBNTH3zEoPpfc
y+mAkRPW28X3pQ//z1tGWj+DFckp0PUqPkVjyM0HqeZEqZHu0XrAbkXP2vKQ70TLLEoH4h/wusMj
t/NrDnPTsMb+MmHvU8yLhtcBYTHta4U4Kth7ku9Ms2BzSQQh16Q2gM2NxrMNEHW6ytnmShjAUHOi
10gw12WOTdX4rCFdLi8c8cFloMWgy7NErMs15BOrJgV9VWJPyPBsDcYsRKURvqQrsjCI3rp3VW5A
bRGgE7IWnnT/SW8EIZlGLV28e8nkSOSl4TORuhIrjkBP57jLMIJGhmPccf1Be3bIgy/+8rNe+F5u
IO15yu2k2ZPo9Lvyp4x633Po4whStUN76Km9TzzHHHLS7WvTZs/tfe2Ef/W5NS6NTQCoCXjP8O/Z
pim6WqQrDNk65S0+/mtU4zUobda/plndWsGEl/p1Uj0B5AZLeVNGxKjMdZa9R90fb4n5NdEjlJmY
Ow5i2iEdGy58pMdbPrlOj5S76l2vvqXqiK9FLAz66H1INnjPnSWtjnWHCeXgmatPjFe4JBXkiICh
hBbBhmrVzlsD4GRINQ4z96K3cvm6Rc5+Ke0H1qtzzZTmPdbaOKa65IliVHBK2B8PADOqwPKg0rjG
OfN8YrLgDmjyLXlcFIOG1972ptNveGKxoFDx8VpyXuUwg8uDPwAYO0Srq6nFjfjT2zIcj5bAHm+x
yw40hDsqUFWJDcfYPgtiRNFA6mCDL4c+ajmKSbLlQpwqjaFOJ7RS+f/bn9imBATs+tRYgPoLNTdI
CE1ahGwlh9s83RDmrRmS7aSRFkiK1oQn775tFOydRq+ZcmR945GyOyQxYaTLdIHPODbU2iLIrkHh
PbCnsUP9DIdx2cBisYPFUuw+jESqKQ+iF15SiwTz/sazphaRnsdvUmH4C2Zea9A+mgNbiLjdumV1
T7bhiwOhPsr0StivZVs1+aSqnGQOcu/WnlDbLg/W4ocX1rxnrQS3izEAIAPMN/Kklk26k+bCM5D1
KekuW8EhHAnUmWENoCi0XiIWE7m53mnKKuFrraTbA8/aQyVABkQDeyCx6q1XWE/flLVCDY3L94e6
TNMeHeCF+1kE1Z2yyMEXTSzIMV0ZsI3atgGOgX9RyZG8Cf0GPqE/QVFPrteFknlp5iYnePrPhT2D
IBJL/yUeU7dZCIWtHJ6RAO6VPSNpyOPV1BDj5tmiQk/crUJ+JNhqaZmSmN0Yv/KQZa98fzDOctcH
n77UiBTlBZs0tJi9psKGF7XhJDQuiLznQWezVJdhywHF7U96dpU6dcgLzOzofYqViw00VdXo9xSM
uGLli1lxK9xZeaEnNFhc3yFJNS5Yh8DzmW1z32bnU3KgPAuq1FPNRBVmJtj5g/kFMVII0d6e5YUW
ucid9u+eZyFIvYZ6dr3x6Hi1BMopQX4NRu+tUlADENAhLkBZSpvhiT5GX51+u54ynzdEA59CmQTL
JuzEELGyzoJJgBGVruAshuIW6jHOvqV6wD45rualo1Djp6Xmnb9+VoeqDbcIITmip5VHxaFDGHx9
7+AgxZLREM2IeSj7DeBpsb0aO9RlVFzq5/3QzQNLR2H5SO1czsrVqeFc9pZ8UgAq8jGuvIsM8vCp
+e8MM2DLl52X/wcfYCu/b2+4tEkZBAp7iR5DT+31RhntDzpzWEtxsz9mlfcD9isgdEulx/++3epK
uJLLmGyfFc7tgh6m3nQs8DnAC1J2sEZ0vAgR2UYXj4YYoNuCSvvbCbAxy6XU4kth2zzpmKQqX69Q
qGj5P6x2ZtgL5JhPjv6gRNS+AJIJ3ZqXPXnaLanv7M7Msa18u5owS1fN0FQ0Ubt2SF8Z2tzw4ign
udojsVxZmGL/WxQGUV5nc4ExUhAEZvPeXoRjR5riAwib1cCR1+judtbSwHp2I5Wl+ItIWVEwKoLI
aHB2gwwyN3Hgl5nZ4Lke0d+4AdgZB+b6Dx2/12/TEsCbF2643O0FJPeAcB7YHLmYzdBiYxcJ7u72
5jhsECp4Q3jEEE4ichVunO1AKn3WbTNUo0tR72V58DdeqHBWDvH4Y+4A7l7p0lmc6JElz3jUcckZ
YU8wkbKqBIhalxPL9tm6bmkQajlIoILGQ82hpEwBvWOeoCi5tyRu2VrvlF+WnZLPnp363X7kgwGt
ABxL8V22KMUudqzPREBzC3XzklyKR4vWSlxJUFCUhl1x7kfIKjXdydA809WtLqiyO5urrhvp7ujc
6B7diQMjlU1TKxs7DhFsNwfF9WgVSamSy8mi/pYyDlHvk5BnUmnbaOTorUtVMCNKqEssK5bJlz1K
JHT+2kZadam+rJFAt6ISxAdULASHPFbAdGPN7QxdawZW92zo7jnTlDQFLg/Cx4yAp2A+O0PsQArJ
L2afS97xJ+QboQtooCKe91/s7xWlNKcAfMdAggnX77FAMJswFZ9pi9ZxXaDVa7xFwcN+oCV424Xu
WKwUMNpgtq4OqaRX4H+V44Vp/MTP48itsZdKHhZzj27nRFkhx2zxSkBp6QAopF8EBUSeo94FkdnV
w1EE4weDqFc+cGdqzehyR6JZi0aThcJce0y7/1ju7DRxKbkpIzMrX7IrkmHA7uUAePPK1NvMPNVx
iOYAxrjF93dNzUw/o7oXQ8BG0kxraK9rZhnfeM9fD4ARb9rTdXzgRvwnMg/udk4vnkR81rfFPooN
3NGKlqkbiQyl0c4sGBgIB4TeIxHRwagNiSgu56XxBb/4XUocS73GXQHb1rQ1gDliVzjpYMWAZ/31
J8aaf3EXW2TU1SBMeYPRkpx4Ys0F4gFAmPU3/10KGQMn8gFVH8tEAkIGNsdb8rHiuSORdUxqZ/n5
DzeRveroXjqrkTAOiewtD+B4W4HheU4DvBcLMEbwLp3eRcdVqpkTLKNOy2u6eA8YmUm0JwGPWgC0
TqyI9E7J5IM20H+9N3pTEJTNkwYz3oxTHpHee5LJVyd8O1Zw/PzWRQsGA4bFnjoi+3TFMDVsNFk5
p8fSEFLBvQ6x0CD+XHPmTCzxbykNqQW7yHEJfa5N2FavRU+Z+rjb7CeolKxIRPrk0ro05CEd3S2n
j0yB8TZTdVP0Oen2b2sHAol29FVdbCUab9y5NpYwTzn6HfL+jbqsK5bejIGZioxymyg99qSIeMnV
VoHqYtvVyMc1lcI4WMBwOfz3OqLqK7GJ77MXLeSiu1RdDOvr/GQxgyXqDgDS2aqt36ZtIGZh+seH
76iMb7Rm1boWRKa7z6ad6qh42exSWOCjnSV2W4AYtMQR/gSx8Z0jrP3tbK0xFr72PCr6j/x58YOi
ZC7p0s9Pe3jA0P31w1qWBXABcDCpb3D/YRsY5SVrAiT2bIhi0NKaZiRqBvyCMYeR5/0iP1qoWzZ1
iKvKPmCOB9IyUFu+1W9h/Lhh6qGXxyezSB19MJheJFXT36fcXfS3IYV2EpSV4FQ65hg61S2P075H
emapVb+zxMB/iiz6Jxzs+EEcyWtFa2sk7GEuuMQbM3J3JSgKwU59KbHRfQ6q2bmPzHcFt3Q/qayj
0JCFJpkOIPyKud1sREiKwPFN3/YuYXEDxBEVAWWNUE2juGaOaIBoZSyP63XKw0xqq4enrv/u2FEW
kJlIe3YUekBd+SH3qL3PEXThhdZplr3y6JmujkMkjrdB+E71eYPcXxS51Wao30pDU0Rnic2TRbHP
gCZ42/iVWmz4hV5B6kEqmv5XNITLpwrh6QJUKlyx1TBrdap1CNMhxRT9wMnEB52/xM8xZkz1rgdl
kSMNe6Dzkqig4w/AazkWXmFcdGEjIryBpK3b6Ix8G4nxO8LUoQMPUZQKRQrGwkkgGKhj6jWE0IF0
JZN554STrV4nVgOXe0RWYXIue/iJwdf7NxDSi/RhG6Z0TVmM2f+Gwc27h/q1EJ6PNO8hlR6JEBN8
xoR+CmbV6fskYS/6hK0LXSanwDwMYAxkAOZZNNdlBHLOH4soRIfhUbA/3T6znAg+/oZer+ySv9BG
GcAu0pS4vbC5wdrZ20AF735lUn2VZECDIrYBZ6P/Nah5rOCzN2ySRhBbXcwbuT1c2+7iOUxShKl6
X3TonvGvxXRobtzUBRRl2vR/6r6htM6DDA0BM/o0C5R99LO+8VUhKmmSXIWxo9TLazglrls6FwaQ
ncBe1IGZaJ24TYyXNtovka075T9lJUgMcunzAYfMDuBiJZT1YjMETm9pkvcOudq43JCODFCgxZ8A
3DzsEkDLD81RpCHG+0AcGtFfUILXtSBkDah/EZ2aPrguPHfuxbuj4Tgvgl9yB1fcvwp5SNxejFVR
iCPntJvedqVB+9kXOWK0bSM5MV5w5372a8kvl1KpqXw70lXt3VcWbh1uqzs1FtgBW+aIxjqvEHO0
jc1pM5HIroAfrJbLIlbwApX4XuEw8YMpV0Dfv1CPCfKYRC81F1szEONQloXvF7LsD08gtD0erhtB
SIHkW/UBj0dRbkhbT3A9MyWSZMbBOJMjrK+h5CyDdUlZtbSzHeYr7pHXhpabn9G4B1lzOoQRhOTk
8BXU0Ed26nciujhVGJlPQUkYIcQ6v2+R9MsTjqxjKVftIidJG34bTzQSgdvLxc5aYW4mIBsKzqT6
oJrh8NPzbEkoPly/+67vnictfM4WKHqv/YCEBwfZzrWNjwu5+rqb52i5sstDhBtsL34wx3C9G35z
ZUPmelmypHwrbO44XdJyiiMMVQurJ/C4oSVw25ROTqt9Nib8enThxJRBjosNw95vCLRSrVPrfLaN
8zsM5UD/XbDzROoAhBXrS+kjNWhzALAstbFBvg1AQL0sfYeZSAT3IThKyASQvZWECJ7FavJMQhz6
DIcpp1oNEDe7Eh7MRtIMS/94jy+iQSW1/dh5apyjAtbT0GuZSllhLD0/5534HH6zCoBQJwy0SQku
WurR5QkRQp+LcK97ukg3FVTkMRKjzRTAgE/eHV/8Z/OfgAsh4rVBx1003GOTg4Dv8CpKkbhXCXms
+87Tm7A9FW7+Taf/b1KC/71V9PhDc0pnRo1yZ/BRKrYii4WEh76A8aNzqZDcqR6LiRHuiZT5rmKs
J5fPWPQgUBfPREnCw8XN9bDtUH1mo1wzsM7SlJRAyXhIeP9P33ZpkoYJRMnvbcQs1wLQKcbiE8ou
t84SrCoFzT4H0JFMu3moVUmIA1wPblJdpBiOz5oVpeOl3MAaSrfCSl88x4EKHMVkbw5+myKu9HXf
/HIJEtOwR031B9MyRsun61xkB4yQRrjs/m5301n+aoyZHHO+UzKbn6neuOSeF6M+qENlVrD8994E
7PaLhd4+F8eTnEFBx3rYrHAfeuVf4HgV6Xv97JmSHgjQ/pVgoD7ldb6P3pxmxon3TN0qt/lWg9y9
CKRjFP+v+RdX3AJm31cGET4Se7lRZigMSq2rIpq8Nl/E3lUBmAD3u4I9OyvFMhX7ize1oDLyLbGV
3VpsxUyyJ7RWW23QpqhBabS6BlGNUceWhyfIHatKxX5P6pXGoblW46YyvpFIJHeYYFp2GNzvH+nU
FMXGNXkO5JTQbNzUdGxfJ4E40xDnoATuD7N0Gsl3z136NJsEdDE3pkKwYRXWE85y0KiOIw4Motrw
aJCb2wNAPnRhJ1bzmUYaDRIJQHKqxFF1FdlTiys4Oc/G2dwpoHBn+QRP6yIwomnWkbOLPyy5LqEb
GDag+XbXqTa8cLuffX86mulrSg34XfePnCTWGCUhC3ENGAHfu4B5++XejSu0/lygGup5YCglCTOv
7HZisIUMogawhMztoCikWZfvkBr8Hayg4Eqa/s4g4/xiLmT30rCabObH4stcwm8aGOnUYtpKSTNm
wYg2FYYcTdoBP0KsekkzkyLMZM9Ud4Muf0ipsjgUZOghogNGofQpnRtKzQERsXl/2WP/NT2vfoJU
QNuujuh+jRGzE45s9VluXrtdSkCZpWtVdUC4JwuDAKdx+YcVPd02AyW/mzgnDi1l+4XuascpsvmG
XjN8TWYxec7c80dDDKBxM78i0fScYxnI90fEQgHaNN9umzabr2VdAKCC6bexGKok5MekDsnMfZet
eNG9+puP5exsGDT6CEUA5up+XV16J4rFO9MX66jT8v4JvPuXghi+B+q/XYAOO4QUktM2VOds+upG
ug+UCMiMRJrzCaFTeJVhVoC4mqIOtIEWR9/cLA920G9YjPxHlhDbDZ0d/C4qxzD1FufkE0fFZKFS
EX06vilqL5GIXce99v9Dd0NjQrVfWNqZU6c0u9uLcaHH/DsFjasswI/4YKSda4xD0+QarWjJQJNT
PNNK5hWoui24/5a+vz2x62Hv7YtOUuZtx6uFFTaULDllq/wW9G4+xsgNBUfGbLOCifVYBmi23s/v
AI6gBLU2n+mogMa07fU8R0PpINThcPyTN6nSDuwqKOKKxALtBiQrJcX7Ayx+DEB0Uig3ilIUTKYo
8LHFLWw1NVPM+xHx3BWlgjy9KL6Cj8wWox0K3kAxZruwssEC8Fs2F6VdRe2FlxN8G8cr1yvY5z2o
yg9uUh4gPJFMNDhmZI2Wm3k3v6E8JunM+oizNXh9+1NlH4T0hw7yS6J6fc78EPXoipOlp3mt8fdy
z+O8QmNBBuHKDUV3W0zQJgJjQSXKY8h+M7DzQUrnKq90dkJ5M25WQs45GCPx32jx1bsmH9dfmsuU
QKx0r7XemXzMRI8ZIw0aCr7iTXfBk9mKZOKa2z3uXHZVjrrfY/gKOjuOsOEQ5kDNiVKUckc2cCbB
utG4X2X3hMeEvutiE4aB8p8+qzI2xPxcd/P57yXtes17rSapGVV8rx0LT0KR7pM5jqIga2oOewO7
oq6gapTMTmqvxnedg7nkxlyXDd/8Vz2P2JdlpOTszs4ceepFxAeFcZ8XRGlXRgksx6wwhhresBQh
5cyl9uu4yf/t/Q9106xy4HEMxAjp+A9U285fkRELlnECb+fmiSsHFzAKeIJUaHi/FvIQh4PxZWao
4rFxMlJUMkfvNP8EerslBL5oc75CdVFe9YhzOymkcxrKzWuP5Baqaexa5oYaaqiw9elvbTx2eLWb
LXPmfWkNuUx9pwfNDy9mmXOohIrOVCAit6oixvQLfBA+l4rOdeS+F5c/OZn3rSVw7JLs0nx8d6DY
Iam6HcsVI8fpoTN7GFV2eLmTGN8TdOeshxtoNfdSQApmDyUSobeEBqSAJI4GWWAH+Sid1439ZCaa
iU1bnxlz/L+z27EMQOsgR7Vn+FwQVC3PxWtUtmhELBMRPCMyb9KZ8l93gxoUcuG8dFQ5vXhgJ2m6
iZgzejBpb3/4aW39rHhMW/60io1qxntg9TRycJpXxz3u1sjoHG7YvJkNrWVuG5Y2MSmoVabTzkCx
t4lSXjjNifm6/4p3tVAepZeJ0JQ35I+4j5+J4xya33WW7gF5WKcgdSD/EI5CEFyQ4PmCQ60x5o9H
8zYRmoA6HxYZEK0LFNUVMVrCo/rp8zieEBxaG9UmqPKQccIcgfCCJmsAWMQgRnhdnhwQY5Qh/51E
aaHlU8JPSjNlBtCu6i/S8ewp3+0RqhM9dfg5DTpnyzFILgzomZlD0OSmIx4kP1LCT5k/9nB+TDjI
FGRFMHafBDFtmBfpJnDkldI9+98c/LyaW6FqDeKU74TJzNb+B2/thI70lERa3ymu2GS1+Zxf4mNS
bw9oha2WBqeLPUZwjVNGZtgRiV/sEZ2PtcTZDUHkjmn9zlYZI+xArJ9r/wuhjgqWXSdLaCstlRd1
QIAYMp9CzDYXmlKpV6Bhn8h3isO/rM5NKNnwa3vo3cDTO6P7I30Ty3BmWVkVT/dyGm43PsqaGJpZ
oTrFuxAOTN+vB1lhJ3yg3zaNPMsTrfbV9WY5S3H8xvXzh9aWM05AJMBc0fHW6JP0+QVw6B0+2AoK
GfRhqjW4eFsSNvqlCkxim9HVFSBGDCkDjAF1qHt2DWZsiAuB4sVTWEZR3/klFaX5EXZKh9+yWg3n
UbRP3E7avzmn5s5a6Ct89rbFAuMt2QWInq3RnA/OiQ/lLIEVPz2ymn1BkWJfQSjNof+0lJXLqps2
30vS5AzL4WFk3p4YkIwCqkGR1j7E6aPljMG3xHkqwwegMjPjQ5JzmEuFcXqtQcDr2/5ausEfNAfE
kJtgD0nJhWo6FHTbBh5gLik3Qf8Fdr+GWoZxY8CXrcDS1DvBr27PWaN8hPPL5geLxUfGCb4GmVAP
ClWFkosyJfJMbMShRDJWUQsqJzzG4FpOchy1Tzds8p8I6yATS2vD/VoIINmTTWgSEHb1a4804GDS
IRzS2BmpxmfSlATpKOHvgPsKqZ4DgMO/b97+nz039d2hmMtPg0SCfCkJ9fdaO9yeyD+ZfwaxwmhI
lSvw7WU3RGwULp5T/wkFg2HYV7X7f5YfMzLFzSIXRUMXf3GEbETtQoziebWlPBPqtY+TD3FCqBEW
7FpE8/imsW+ydD5uo91EMNwX9ucDNmxpH0gEaSTyABwPUGIECwvC/TCQLOsZ5z2gLV5CoDKMVb0+
hVK8dJavRXh8Ptsw88zmZ3pKUoxKeyJ1Ynz+mR+Q8xAFCuN/Sl/7qCIdnmpj1Pm/fFNjBtJL2Iry
4XyI1vI4yGfv233N+MCqDnbU6zdjydhKzU5QCqgd6ir6bIYetnqd6V9SFihwAeUgfF/uGGX8mTj7
/kbO/fO3MsM/uSL6Y7RA78p6KGvmhqyuHC1hVzAPeKuCs2ovwvbIIfSpjUpEyxkNtRIohYQbHwsc
Kqm4UIJGSH9xVBQoXw9wHjlQ80guUFyGdlE48ayDfqxXqS32ASO/0jDHrHtKVanTF+46bu+O7XIp
G8lXr055SNNVpB7MhqZiojv1THfywT0X5S4VbNGV0P7hweTrlkq3uenDjUAAMWi4rHkNTmzv+p4l
uELtSqgubWzXQwGlZ+1JYfndHGYwetL8zZbogHNWldaoCYZ/ZtMxsAviBJoUsDU0okncUkSp5Yot
80I84IgngwYahz7gBzx6FGqgwEEUfr22i9TSz96tzm+I99bxOoRduoOKabg2/Rnr/4eLM2FqHscZ
vKgRCb/VQTelJL0AA4A8KSBxfEZZRLR67ISS0dGU60NgvqJca+nX4w4cbPxNlJap7kKnVYpCX+lO
P0pQSt03Ll3VL4jLia7/OcA6OYROdIiEroDYpLBM+w1Ra7PWFtYzC0sgPw0xaxrWrBFBVsQN2X+l
Kq+QP84tlSWtt5gvRTd1H8T3PY4oW9IjOoAucVqa3z3Pcm8ZU6pAidqbwOSv113/GfJ1CdJ1OVCb
VjsRemJD+Xh/QlnCGC9nJVgwl0C6Wz3ZVhusY2pGLJp4MM4tGHcrBNGlYeL3crLVARS0yYwrt+dj
YF8BbPrPTa3p+ZTl+NYI7dLr7Ytx2rXiVMTuINuTNxeJC1kCW/Ouelf8/FXl2rFCEkvLE7RnIvYO
4ltWMBTAMln+WrkH1StQARL102X5VM3dUJ0XQCWAxyoXZGrwElf/VTxllgqEJJkFD+5K1jL4RLF8
/PedpWSTrrw+mdEDnRNtVlrVDBgScBIah02y6Rf7h6XP1lGK2T78htN1aRRWLbcYxtbjM+Tzy/2V
Zi1X4Om4jfeOKHKnIw5gsNbC0h5wPsvz9HFXfYgN3j1lMgvKNXmoPpBFRxQqLSWyihmHKXlkJAJX
qjUL7eflAL8Zt2CyGnqiRBfs/xlxpcnCZYCTppLbGhQkthWZDOm+oWMir9xe5kfZiQXtYRoNDcXl
jqUTNr7rNNb3phS9dWJGRtbz5LRhYdde55/AmA+GxLONRtpwpcp/DjMQC73CiW/BzpRXW5zGttgt
llMcqsqA1zk9YNcJLTlwtibkccyGP90IovMW46lbuz19+6jAwQfY7CyvqfTIl0/eg/XokjHw8lZI
d+4NDN1uEPBmL//IAu6ik365SEoOoiYZyjXRLVa1Bf6wefIYfl4FZnu5mgVHzFR4CvLgjReJmY5b
0whXLNzducE6C59boE1aIEOJ2HGQSjsQXL1st1ReI0ljrnaZ/ysu9jduxiaVDHvJpH/o8mhUARFO
BpCaYlS3xhRUmQFmjaXcVhSYeZXhI8puxd4vluU2P1PJCZoW+MeRhSjmmteZ9yqEEgB67rLkTDzH
NqM3IaAkHINi7QHHZlJvOubRLotsmqUQ3w0VRDpmg3wzD2I6fWyjmaomO/HIKy8wYySndxunPU78
OEuGzHDxhStvAtM5aa8qjnWAiRWyYTy/AjYeBLMuTG1gnzbiUZmRjmHnKgoEjnXUwfn/gw/SuZJP
YkyGnCMKUj24PJOKWPUbigRhu5RFM6z9eJ7bRRjrTvAyp7ilqZyIYavyG0GYe3hGXrtmh58we1W+
edy/AFhZ9j6z9QPsOJ0em5df3et7b4V4LK5koamqFc7mxKu9B6NHi5PbBoY6zhoSF1+Cf/qAMpRJ
mbkdpkc4FGcwlCNzXNPTGTAaiyTrJzMw2WEoJknJRH7V6czgMcc8wHA3ZSkpZq4RgsznnzT+riCD
7w2sY7bQx1YHXFRFTnEtVqWmEw+e5xIG1ny9XgKpwy5Gt6j4i7X9KROIgitdBoUo2s78Cj5t196K
CvSREK4ipGWshu4+LEnv1bZxrowwOXgafgIRMc51QBj5gocfOkk37V7c/VnMjKdkVYXrc26js0mz
japX71EDkEl/rbAcxeOirhwQzEFw0tqEVqLQDeYgXkSZyTfyyg+eJJIzI+LIGjkZpyzsuw/I34zM
7lcacpB/ezfflIFT8sBOs+bzAsOoy7Vt94LaeLCPHCsD1whP8jrcohC8RO04DXJpTNuaCUkCAUFB
bY3vZefF/vx/HFPTEJYPpm0uRWQInsR2Tj+ufTBlZP+NQXwmBsjj8FICtWnGgv4j30lns+HM/wgj
9EHfZhmayQyG5O61d6SnHfO6nuQas3uQxJJuDfbzgvkyPCWvd6uYUixguKFdN0fNNGtnAAl00BV1
AGEFdr7d6DC/g6QSR94NpaRmIuiMRnhBPFMEO/GJuPpndmlJ2KxRMvf4nxijSdF/MD2gS116CYo0
L010fCyM4z9PbzsBlJbyggz0xTQCyXt6UBDE52W1m7Q2ujkMx/YibGsv2cP4jVSv+AyBndqUtDSV
4dMmTFgIv9b7tDtMP+1eFXsl4HNYvjhg0jioNXWDWA8hbQLuIGcnZ1QErDdFF5EbIEn/yhhfK2JP
4xKoYAyXnb3mNwYfMsRjpxwiu4HMwDeLotyhTxwfNRs1nzuAnSQL6QNPQD0qSOCrFBqT/Gz9DrIF
zxQF8HjSoRnK5JF9eZQtIjjpyUu70OHKQHF+5+A/CbCiAABKdI+v3YVN+jUrOEzUmAVki2C9c7mW
BN2ZrftCtjp7IAVPu2PIVu8E7PS4lG1k7VbCuVeGMdAYxm0yEnlFAfvA8G9CLBh6ZjmhPhttq6wI
hAy/NXpgV/YcQFTdgwqhcWhkN+sRgZBUzDwLgvLMmnl/Adef6ZODuM78OhBooMX9Ud7DHhHPYJ0w
WwjtkZRe+U50x0gHVTSanv9bNIdflLWYssQbfkdk+LMZ1AX3KY/Usr5dNFdWYmWCUzZlcpRSRO08
ISykus8Vq5nMTCYyx4Vuckzjv/vjtegXe9gwtI1b4qVHN1Erawsz/aqHUMVB9jVp2l/rho591Cvu
PmBmKw2ZLqAKEgOAH/RwrZpPoERC7a0AiEA+FznPV4eLHWN33HVmceFFRFbcruJGnBRwukbLlkK5
yONpVmmnrxI1Qc77IOJ+42kaXT8OpXEyq4WjPpn6SLuyJ5hiTeYR8BsQSBvsWSDvPM9mqGgK1OZT
a4Ibet79h4AUy5UI3cSavQD8IYbnYlJlY18DnVeaa3T3SAka+Q3tCWpN2UpyovH4DvoTWUZsVSOt
DSRH4YKry6XUJdtJpgdsA5AZIVd244tx7jOi+PIpKWgkxqG2q7vOwvzqPkZiKaYKk7hrHCQj67fr
PwUiBobhBc1xrXBDWcYUOSqMCcYP/Q8nmxIBmvMyXCRmn7AlxeFE1h872gcN6fQ6RIEa/NORUCug
dmerScf9n7c515gwZzSqOozaxChntNtweARd2NwOFTfZ0DSWPP9ZaS2dym1xBjg4nXBCKm6SBOon
0isv4gX5njXNOoPT5i8MwCpH2XEgMdnc1caJdM0VmyoQ+76BDS7QxSkO5sXqQ6VJvHxjINk/j/VH
aauG16oGqkzTQ10ms14YgbwBiCNqjaxCfTHw7cwMA/znxnNUC9bPhlEhfKGN3ZdJ89EVY4o6FBM9
YL3zLg1xBik/4fjAT+e4uVHvvNpUcWqPOH1ttyfhfe93ujbFyCMgP/Ey2u2/omPmYuB2uNKp/neb
gx6qgWEcsxrse6pUYxTML8+JT2j6526XSsfVN3OOAvSG5oPgsg6xExUdz1jDgiznAv82Wx7sTnrK
tY7aonvus0+eLbCXEod5LFyq7XWUA1noBwg2DP515MQdFAxjpRY5pFvzHb+Vyiff1OTKuB7+VWjQ
YIuO6Ap8bUpTbGjcN0kRj4BuDZL42GHVbX0vdKmQgrF+FPxL6ZQZ58ua4dS4JOxzJdHG+/+nrT66
mNqxIzpEOYgZFYJVAaN9mC9MSDVfoyG/mtCfjXaIL3+dwqjjFmXyq3RRQwxnnB0tU2WDZKeviC7U
t06q6TyAg7A50tYzrpmnpoZRHvNnYPLwvqyvvmC6W0S93Loxwkdsjy+1KyhcUiM0zpaFHkiNU/Eo
fjrYPQCK2vCe4Ju30fd15o96+UE5b7M6WnqGEd9XhMWaYkXbCUgHfgAlaShRn34thxIAid+nBk3L
wqapt6A9QnBrNfSDgXIGGcMJ2wruyWHyEpsSiqO0ureiHfxAH+qwXozMwe+dOsFlVbgjaaDoeyb+
1QOguBOhsD/Z9XI82pPEUyz66hyktcfo63+px7wBC4d3E1lueBakxxjMssFW+al7c6nF48kb4NTZ
U4WDBu/NWe0Hns0JJDMKNV6B4VX+sV8O3dpnRm+AqMD6/v1FdGxmhG/z0CftyEhkRH25dUOP6tES
w+tmYODFUceUt+OpkVSyG/nrUfukC4Cd7xeKt6NFGvOhYt7v84adi93LUBfIWETAvraHfSRg1h/i
N9y/8O8QO5igdkXE6S4fLhOBiRkkH4seDWenN9+0+rJ8FKzcv7jktEVhO0r73uH8BcAysEJ5s4aZ
B6rG88ZeiVkvg6qmqeXgcX/P8jSWHCqy6Kl6elJ3QzWFu+MXDdQD2xfD4xChjrcrJn7sBGW5o4Ph
cRMrANHvLtR1QJn+M6x2/qIC4o3AVCwbD2uq1s3nGPRajkADor/qn9X677XmRuTE33BohTbyZ7KQ
iWKKj33r9XW7sLmO0yjOBDk7/zRgCEVWc+gpCCAbNC3EOFh8hqnTSP7sMzxTrb0Dff89FdKSx6gT
8uE3lbcptQXh7JsC6YCNmF6NZvc8s9kPmfzejVhBvCYerGO8oCPa4B9fM0FopVcgmQ9V3eIeGpCO
pgVjeFcD8Whk3juKPcfphrAF/h6q0qHSSRRBhEmhWJfPvy+TsETFlyB5B0tAps+fxKOGyyekj8NY
/41vm1MRmGteaKao36Wg/s0kTZB+WslVEn46HHPMDHrsUkxJrsdDs3ZwyU57bYia8YEFIKo1+lkJ
MFImuK8Fab90HDhco9K0gMkPPF19TiuCDooWvo/LXxBDrQtlQXv1Gh7D1qJ9amIKUOWAExIrYnGN
Eigx7Blu5c0syqWItXDza7qKknAbPPPUGuZLSb+pidQUK82hGatXwo8LgGSdeyQ+nucL8COhwhBC
mmgrKXfvye4oMOBbvEgSpxETapPZDPaNpBsfr6aW/VBuxWouPnUo0zbyxCwcWyJoNORNRI0lRByg
6R07Jsz4tLbF18CrHzvQTtkcANytpBlPO3ikPmk5NT8XdJ/vrFzhh8Rr3qkIahpriVKbsfYH+Xyh
v2+o99RUE1ZBstzHaAn2z3yOIyagtyKFoOw5f05FpLBzuv+6b2ZNz/sjcCC19IxsYYoJoWGdenhm
UjpCd6n6zJxA5dGtE19n7DQX2sCB8qT+aYe+gNVu3/lbkzzEzKrKZCW+T6CTvVrsaS1eoDiin3yU
3nNoSoSnOKSPCXknqT/L7H6DJFl4cXiAG3JGWjsz9MKHx9txEfezYmIfGRhwnS0DdCf4V4jEQV9S
x8D4RzDYIAcsNbV4U+e8MAvTefX7lBiHxIy3dbK4iC/hb0z6qm86p8FFw7EBIc8EIeyzFWqcTyEd
3u/LiYTOTWEbHJvPZVd4ABFV+If38hXVfhUPoMVTaqc9/gzsAlTJStNTYYzXEMJO/8m9Ezs/R+5k
KJaXDRHyyYHgn6Wr1cY1Eqbtv/K36qOUQBoB6wZoqwerlgJZtautjFfdOLYLeato0gWPq1i/L5+y
HYoV2i11sN9ixyM3Ls+z/oRqhHNHgk+KB8s8hGJ0goyM643OAjhgOCOUOQEuMMqLLkJw6MVxQFan
OeaxbO208zorCr3ai1Qf98zKtvMMi9m6X4cRHAyGRR8NomJs+6GcHnqd4hKZgXxu5O6Har74QwE4
fqZpbaOwLnn/f9HLT6LXjLNeU7UAnlmkrNj/DDL4qS8s1p+9XrZj8CZydEbLkK0KYPexPci1UXJW
usxK8v9mhemYX+M6zMLYYgRkfF/boKmppFDzdTOcsq0s4FQgVwhiCaWcQ6ThmCR4lOqG0kyjj65h
FHbWpckVDxuQwcyeTPUtcd9qnY9DrI0j8oPWA8iqVzmsqsBv/2Wi+JQvnFXKmrOAjhYKdnoXqB+5
wMRD+6oxyQNmF1m/FI4hlbODl20QhiCbEL0YUEJuodAndRRH20VRGkev+HvaQaKYV14bvq2DzCV9
ClP2xuAsuSm9fpSpvkfhlo7qRPP9OXMEUoIj3aoZZlyOgFm7clF+MuEk+SVk/RTW+AS+/Yk2f8Ky
ssaRwIxO2v2Y0UGLFHwyMlOGLvSs7yXDlKvBxVEqduxmj/JECPTwu8ji6jXCDsATeZ6EgnU9fRIr
08jxyEssFP6xR9cYUAUuxa9bf8qsDJXbX1OIi5n2u/Vly3Y6JAncC/yQEGqVfbpBgg2Ycw1dmddc
3ii83zIQct60N+1GN17zlVXllfSsrhdDlQLE9iQdoo7/lv2wIGwGSlwFLqfgvwGHS/q8Ef9AhRyj
+AQ5Y7T72CgwmepJHGQzN5NsOF+nQahHoMbRGh7Xx3mudwE3X2rjYaD/RlpbWnszej1iS/41PIwG
q5tMgW0dgrHCCXfBZNmkNaE4kpsbSNA02/8eSPqXnkY+eHVR8hN6/qhpSpF76e1vYKCL3KUAFg3z
0hYNxpA0a9eIfIq3hDanKdeKjnmOBkcILtmG2wlRUOJ83Z2jK8x+cnZT0hnj2cNMhzfYjBC74FyI
OEa4FGaZIiy6/Csz2G3MDMrodAr8Qo3x/RtZ8tkdnwOI0biZ8gtVkfBMKep1m7HmpnstLaPzlmzU
DK0XjIz9fqLTPbOdSxRiHJKQMBaykkMvES2eDzwQx1gRBkEwkO2SGNrEVFHLdi7JFl4ddW2GOUnD
xpZfzVYiDim2Z/5nyg/AKJbI+cEQftrLQCbMzFcLIps9QPjw+2Y4xfHDsZ28CkWZFH1RqzmtMQxk
5dmfQk4q1PmlwGhwzHHw72mcCGQr6FF1oK/XSuwH4rLGIq2zdMdjQsjGSU+YbNHi6S2sMUcl2n+4
GMnXzwH3/9hZjJAHU2wS7L0+OSDUTtGb2U1VSxY05aSarRgtVgUH/jcuNVGIe8heArojg4dofJ21
QHeubWeiWmPjhWBn4q8Bzp+Wq0CW4XSaQoV7r2Bi6aeXYRfwdRBUMmHZqwMsZG4Us55YlX+IAi8T
LTTva0IzDExjWmFEk5W9AnO06DPAqM1FTMny/+yEBnQpVSQ6c8oCw2ckV8Zl4MnLX41B0Xg/HrPV
q5yVxdpMKBtqToJYq8++9as9bTABSNEEOBCO9T8LZ03p1H22Ph/6WQbdXiu/09FGrCJVMq38D8Pk
OTm0KYTdzOLus2y/7pQ02XoAAZU5UMf6gVjXiNWxx3xuvEuTdWPFvyxgxljsVe2xeg/4R456NP/7
BzJuahHUQfOydJyK+l+2B0akMcc5I7IiVA5OG5bs7Y9t/alWVDw82XNMlsms1YEfeJdKZRfZe3iD
6Z2naoEej7Gf38/OcisfjMax0/RdiGR4Z0mH3Gnlzn8t3H3/glpTvaYUemiHWUJU2IlR9jISkn2L
LPiXtP52X9AqngL9NP/1DZ24ABO4i698z4kC7NVXiEP5oXf6+0W3fucEVVg+zpLlWzEm19H/kMNb
9LXalZ+pYosT+/eOHgd+NYW02vyMve4Sio4n52P+piGWz+0bVzXv/4bqSahXZxghko2VMTZU5UGJ
w5cSkb5PmhOGwvA/5X/FXu1AefhCzd5OhJhBiHqnCgPI+MzaLpGKC68exDCc7SC0Hb+KeVgizsvC
t7dnl3Tk3jPEuTjBp+LEw2z64ozEbOr9+8xYdOvB4hZu/+sJyexwG9bjxFjBgwHIzDEXmi81WPuk
NW7b2MzPsgPZdkdcsInKzo6PHQzJqSfis2pWVVYpza0UpouTbtakqlMzcl596Yv58WplBzuNVlYJ
EIHLB2cRoR9SDeQpuhnygwdBaDRA8ns58IJ9TYkpaRpTrO73KHrp5Mfxx9M312SB+hTyXd+CTsxk
0kTKKSpmzwkpJYbjWQ1Towj1mPzc618OMXyHyiO1E8f3fIxcErsMerEqW7TXRo5T3Kvrkg3XybrY
H//i4LjLRch66hUuYeO03K6nl9MCj9CEzNfqXwR9x7nVNx0QqztAUK7XOXfDkTIVnpL5a7O0q/nV
RcYYkqv2t7gCiUlikCwXnGAdVr51job8Z6dsaWMDLL0Q1I29MgkgOZThcP6qOJiO/4Kpqn0DLxO3
gofTV8GJ/ou5yyjy/WfziuOjIOJUosq8HsUv/XFI78QFGZo+3zRZmfmumgUNqjKLsstu1kLv/ovy
Ax2XS/iEpf9AndT/ek327e8Yr4UyECW7YZEsiDYdDCA3dKe6GV2jDlhzD1tcKGviCAy92aZ/I6gy
47pPvjFNG0mkjrG19eBZEQzbApTWP6s6ltYiUsHId/wx1PvYeK+87vxTk8DMr2OgXInbyTT0TNz7
i4inoZ//dSS3f6M1egEt0yVQxoD2TSZ3C2f6OjCLa+RIQ/q2X8jHjuTZ+A0k+t/OLH/Fko/7TXZA
Akxci8efxDtzUIZvTXec+6bYExdbjhZpxg9cZYMtD9UH0jSpfng2+4USN9bytAo8lWIemXBTY1P+
WYNBqtJEIx9zEBBVXbn8EbIKuu9JdJW0HJlOWtLXZ0d0DgfwWj9MCWYULxrZ1cL9f1OXjGDu69vZ
BxNWhUG3/ChxMpNsFXuGB8ekGMoZQ+ljHWoyDYHgGJacqs/F7cqKHgOgDHurs27Md1Dn4mdpK3Fh
3ZduXjrN2eYscnqMByG5S+wAnSubEPrVS13ap3EHUcAQx9mM0zeb0zE03JqXDf5E0lqut+Le4p5t
Yy1w+DadSO9GsAxuWQc2Nq5MuIvw9cxosk9i6g54axwXJ4IhT2F6PbY2UlHG+th6CLq/7ykGskRF
tDHUwpJ7IMzUlnRnAyTrmd+za6SPjGwuxKCll0aj/TQEY9E2h4SZO8HYZcwBxfeigTOk+ZBJWHuU
Y6lx42DNQPk0nLsy2x4K5D3r1nU5g3XyuEBx1aACk8pONABlGpFpYtgknqH8EtpcNIiKRjNHM42w
gQbvHhv3/j2Ykx6Dq4uikcqJs7Olw8/0yxkshmQhoNaiiNxH/6tu8AOB1pw+oyDecK3CHFlpFddP
u2z85xGkAm5m40aRVE5t8JoVeEG8qRbBp+zC2HgY/2ast8CNU5lX3ani3CGoZo3nY5krTH0rm4D9
t+vJs6u5qy/Z2Adn+7A5Gcj7mv8y//+EVV1qPtI7jdabsULXH2gBZ5bt1uyGhIJjbnEWwyiRXIoQ
heXjbkz4IJefncS/dO3/W9PudNasJFqdZVEIx7I7USzJbLDi1NnCUpiOgZuY0zX9hSFBHHsB0s9t
pM0xb39lVPoB+ljjTf2J3f4GDhJZPhl7g7wGwnLmpoZy9l2kQe5WqzqWHmX0tApL05pG4NalstX8
jxCJ1SC1XsY+Xf/5nC7WqBbepczAHbhm8ninqYeovowCkV9J6r4mvHmuos87cVx5Rbtbty3CHfci
TnY6omss3ptKYbvpRkdRTG8mvqKEO5yW2X+hFGDkfjdWIZRSxNmysagbt+bjQFV6z1oQsGWSiR+H
aZB/7CxnJ+C/lRlxVLet81jA+6srGckHdD1NdduTDZggMUwZE8yWXMTDLcnCp27MsAdxhiYi0jw/
6YErwE74icUlK50BHMj9T8Q75eX4ytVD72UUWdge1AjXanBETBExyA6uyEHLQBx+ApuEJGI1476E
+DhhLM0HQ7l5y1MK3RlWTRvvLkuSW6SstNXAMm1aZ5EYPCDAr3qYflkhsbM/YlmeLP46R5/l86uW
w5E0Y0/OL0LHgOM4FN4peOWvnKnVGu9tyAf1qee4zEw9VFciBNZsROwhXrA/Ench2wHNCKCYfhEx
zJwcI6C8o1AxB2uP9HBNB8o+CixMGh/zHgVvbIAxMxd+U5WSJZgipSMjfJtbn8bmf2iE3U1FPc03
zDvC1kp7zSZTOgrzGFxN9oyKOWw8Ps3ChQV9aAK3FVSZHN/RisMiq7VVMTuqLMa0ingkDI1c7cw7
gYgA2lJ6Y2BGEucCqh+69LDtdK0gt2Y466Z9xP4vL35ULeb6JgiRWLYt8uBV8tuRHBj8/gdBxpi0
64mBEiUD1y9EWvhFT42mPJhcfew2pq14uRlVP48VHMIgvca0NvcbELgJ4+hjNVXXZDGDxyaq3ptM
kBmeBcckGVwnvd0wND/WIqjI8/svMOjaNjCM+EdeZjqbmJC6b4Xg0YpsnQB4wNY8aLcM+qmpGD8U
PzdthGIxPHYyFcLYoXNlGGsM6GMb4zYrP4psoZExOq2c5FTD3eTyUYhMxwUkaaVzv5+9nGcg/REr
KUVPw/CzStmAzjTSEzfL1Tcc1O0UnTDAkV1Toi5/gR6A4GTdWSQ2tsn+pWJ0EFhUyMqsawsKxHbw
aVjv4RK3PyqBr5wLFKB0Vf5huV0hOWX5lGhe0Y6ojDjWq72XbONfeH7MaQyW/9Eh8jS35m387GOI
FBxpzlIEF3dBR+nZuMk/qIbWbIQT6T6TXv5B3ifVQLEWR9JeLLkW1wyVw8Tv4eJCwhqxLE4aXOJM
N8mGoM6x6mK3NK9EOmjZAcKKMN1XTXzqgyoBGS0Os8HqwjOdgXCVqt8j99BwVecx5kHyEax6EZqa
kEL9ygmTeU1PJyiFXdvAOpqrp/CV8WK2YCQjYdISTJYf0QOEATU53ryfWUPkBjYXPuNQPEKCh1jz
EJxEwHHBmDqBzXP6mCr/V2/HlnhP5cs7fI4pn+3/kW5Y9cp8Ji8/tuEFASlz+F2zhAyGpBI6qA5E
MXzMZ334RA1kW9Bv+PULEDPf9K+xPHfskQ1WP7nOcMwmpcHAGJszTF2bkaUvnzXDcgaMjzv4UqtA
nOjAHsnlwleWbmkDz+xZnaP7n/X8VR7t38S1ywRvPcJfbPDvbG5ns0Tjw5zPwxeLT40TVSVG60CH
W6iPRtFXgvVQD5UJUaI7OgzvuWE1Inr2KSNe2fH+83hYVTJgLwUrwOTYjC85ikj268VLw3IpBeB6
md2BKwqWloWpVU0soB5Np3bm/cth1dozJzHe9GgkuZ700QVdAdlORIpVf4pVxF+sQB3+ChkIZf7S
os/pNg2RXsPJe4T83kasZ/kHQFFxZdWeumOUictD277KafNgM8ct8XEiSR24iLe9lAbDaz931XZe
OUqUS5X1lNALhrMhvGhaWg6x7QAchS6HztQtVxdHW9/2XOECET1pmOhDIeFWh6jCUI32z8SVT+Zc
j+jQWgDQOlZQrk1rlj9D9lj5nFFNnBdFNHHwSGa1fxSdxKIGjfkXHorl6tvVAT3L8nBUHttF16yC
xjAdak/UeuMFG1P8kRdBvYWhAPigqVBYp/o/JY6XRu+DpCSqGHKWCAL4n1kJpTyXICC5/tKsR211
6nUIxE3to2yCpYYoTCipCqMz0CnM6KwzwjWw3Ka3AFWmrrCJeiu8PhuuPi1/iAXWcSL6fxXdFfhB
W3XsFJZJsNB0njkw2meL3+rl8FbImwLkua3UPys7QKF+rqqT37+SFwNiqMXP/QYOnIsL2jqY9R/l
/K7FzjejPUkUTfLxIceB4h7Xv4YOOOAOuxshCUqfBelCfYaqhHOO+GYSZhShLdN0I5YKEtiq9y3V
inldZF/cta4487E+cezJMdrthzCSSvZzosVK8wFv3uDyG/zrwWAfNRGeOGgB/aVRn5va4TFkMZD5
du39zZtkZtPmjQqHe5qMru+qe3TFuKmSK1wTCBGh35lCFyVnHUa2OV9q+8KCvDT00kl9ZKgo+Wve
MKN5yotKfF9YiBQIWB/XiDUPOhqd+BzaF4FxLuKlJR4SQ316cjTokCi7m4S7lKeF9aHIC7aJtmrM
lgNGIGGI+PN9axd2Q+MAuaZLACOj0rO7LAUxmG5n5VQxeHNXWU31zZnziX34P44b9c6mgji4EAlg
tq6HKvGqUismhsOlWcRUGs101aDMIfof6RLEzj6mltilGj6lqOWbdZvDacgiPzilns844hmLWFM4
GnWEKUded9dDr9fVEeUjtqxeQJTdrfc8C6xYu9heNytXG/ZI3TR/KkloSnbVatf7tcIFTeejVBTG
wXD53KAagfZHtHYAfUdtNRZOFc8Rymi1CKPTs+0G08UF9RfCLtV6Q3YtLOxo072q7U5PC87aF9mA
kdw48nVRguyBSUfdL8I075b8vyM0hLVMlNBpzH1RNZihHZ2k8qbdmlpdbkEMqy8t2stdikAsdP7Z
+sWqBAlNhCWNhRtPj2Z/C9fBt6JgJIuL1PvFp6/N7Mxgcg6XcNIRtql2wiYlQG67lfpUGJ/Hv/ZP
i1molYJIVR8eS5hfMY6OCpwNNXklCBrQokRduZVt1ker82I+t88bzyTZ3D9BnOLP5ms+W6l+xfJV
W0I/JrNtUL/lOzXnMYeBbSFa0t7ohKdvVYPPqJzQjPT5v21LCJeoBz2YT1u2WqQ+qm7ort/MTy6v
UHNwz3W57uqSGOG+ydzep+cx05/zJlgbJ9z/rYwFVX/Lcio6GdErdxJthGnI5TJjzv8WEUeiij4E
xhNcCHqdLd7g0xrRGyE5HoCo0D87pC7Vbm8YFo/dUhbPr4FkJozJLJ9Fk8LjZWlJOCZ4g+9qlJlf
l/tKUt21pBAgr0oZBNr1bP0kQguhSLI8XwmmRvnpf9ae9goPApf08qWmi8YK99FttYwp0ogG4nq9
MwVf97+MYe8aXdk7F6jdV/S7weIyFWK5TpR2wM2X2+Ud8XsZEtxABQ67p09UNfqSuX97uH3IB2tM
J6r2OKuo0TatuNrFe+mL844X9MO1K0Wo3XZwXFMApogpIP12KVSCNuiSIHUBXr27z0SKuWogLFLH
qlQYBaS4X9nhxYjodxcrmZG25BNYelmunM/fQFYPzpAUd3kPCS7QoEObsrlleGFlnkswu7iqUXbj
0Qe5gjWC0BXZp3wvbDpo/4gQPKX9PiGP3Re3hfk4tz/lEm0N+JOp1N0RsfGlUNRM3pkOIZANFthq
bJvMUYrV6aXs8QXJoA7sV8JxUYho1onUw/enbImSNy/ix7PN0bQlzSjIq3S+2lexlkfNCIzYQTRV
8X4tEKrNm5rC8gDY+oHWcr/F2VipU8smrXwZxGtbN6PL7Ovohk80JvvhEmb7XWevusM7vGsuVjYI
bxGK+Pk6VxkERm4nu9mkQFJX4IInT1EofbQuvBXzCrZ1bCTYtx5aGFt0JvZo5ACh+L1hI7+ZGBus
nFGO0Pe+gk5YR1VDWdeTH09dhp8BXc4bHzkOcr2EjAqBVwxvgHzwIACgTTFy+r59WjbKM0VBM+JG
Ly+NtLbL1GtLK4uhJ70gmLaxK0fO1dWw5ANu6Lc5IZtUmBM0LxurUc6UhyzjgbwfPuQ+cdOlL3Hf
sR/T7D1Of1TnsJqDnAqmVVl0lc0jxXai22OjTxksweChDVG0bR7e+JhT1BfvW38287PdB+43dIlI
2tZ6gCGYTd5FbWcBnhrt/0N9IhllJaUlMgbjY3syQPW66eWFWyJZHsG37utx/Ulpggz3XYlqPOJK
w12XYFm0hitIGUEs6/QwKac91fXn14BdIS4agrse+IWobDFBv2r0kL6UNJDXqrmWNpYJ8wPhj1Vh
fX5UtwGHTln3uwL8ZT/mBOz8JbTcDwAm37pK03Q1tApdZEfeW2AwRCzLr6A3Jn2BAUY7rBk2HXH9
qgNSg6RcXwU/umLKjcmwxjSlz1cB7gHMLVRqMHatifwTtWmBV7vqee9w+aPtsyim9IQVcPEFbF5C
07VbYMQSN6MD9E51L0Hb1iWpIFh+q6GUdHrrcvJOfpln8nhNZmokkNrBBaK+CM6BLBnLvmQXblIH
Yvf6QVTG/IXBaOQNXPy8mUvKV7QxoIkrIpCJ4A5glmWbipx/k393b+AMQDvsWawrt6jBRcjps0Nr
kyuQIIZdmgOA1NKRve/j4X7gslEvd90gKiLH3uhC7xNETxlX/KKDqvBqIq8NUnDK4lvrBVwvIuKG
UngYcvQVkhSkVb2QL/rWmNgxbrEuEUkF0RS8Lo4Y2tJBKTTOnALNCAeHokozzzav2UxGm2zdb7dS
4Y554oA6E2BNK88zcWRSolEXE394Dcr2giKHwvmnD+3KwTWRlVfDjyWho+Lsud2keqL7Xkwzfe+d
NXDXJndDIAY7PGCvFfIPWgIfTRn6BBqbguou0yBFIf4BBCmGQ63YtkIBP7PREo1PAZfGMJJy3Cvm
/LqRT9JUGy9zGHvAbwiYUDzpK2hclW+20/65LVs7vCNaEJ0gEVi5IMqEzYmzWjfulR3AP4NxPKIl
RKLdO5dT3MSn2YK7it04usiAjJbRIIP3+iCV9afCtps4oTTC+IR4jgjwDWV84M+FFRFgPutYD4bo
0FfNLf206iq62n62AtQON+/88ml1ltgHISs6G3jcS+HjaO9/a21+HRSwWYHSSnZrThAJYeCqZVWZ
DybI/vSlRUNJCR1kWsH+01qTGbCYGEvzNJvuPcB3OppY7MUAAKUMOV06r+aZAruBjRMkI8umsqqQ
alCw96e8ZnlhIIQEmlPQ9azrhatzF3aCJECfGGOBgsuc/frXT03CR3EgeDMGQm7PA6JYpyvRXM4R
GRF2p7mszN2atqsBLpy1kXnmBNkD6nGz5XLrHbpakM+snvghXfqYQLQAg+RnUkrURhu8c9lY6cD/
3FCoodNfcq2JR667H+J+FT30QKSBW2VTxmOPmJpMyAyn/Q0dYDobLNam3Bv/kcCI4ibChRGHjVwE
VbKDPPHzbIqiXwC1Yq4lyY4SQ3tODoy3z8gQbBvunwjgTu1PzN1J/k90a/zyH7k0zNaqmlI3HIlY
tbfzPwJ3pMJwwsW1OXlx5hAs9PTLjJJ7R3oYNhh1XWluq0roRTV2u+SzvbXgdTeKpfBwipD7y4cT
XYsgo3UorMwSxeET+EvxHX+Bh7mt9L6njFCn1QqEEFha1MojVw/5ezp+qZzGm1p8jR/ugvDKnnCV
3ivUn4B1vgyvTfcQxd9pgYGLI9/ixT9OLrXc4gGABl1xdkqW2+VSE3b+Nf/0CblOpavKrFy0LRYY
cEK/V83XbiacFR/SNJuhwG/x0wrZempRPRh/WtbYm3ST6IcmCFGhoeFuMgFvfYuRes2BCcjM0+A3
ajKKbwoiokImKvkoJZWQI46GLUoyDK3XyxGgmlN/YECSq/XFSlRvt7S30Okfl0l0N4LBfGBBCpak
jOyfGT0oWUOO3swlGhhxzXT85NEAyk3mIRqITKV7W6MXPG3cjh8vU/DbXGzCf/SJamL4RldWLOi2
RqUyOcpyGgX/nS5rNTCkUCym4BOYVi4QJl46/Pgu8yD5CTdz0Egl7sH4zB73rMx8oFhrgqNyBGWh
/uqJaJEqjqjzarMzDcOHt58b6TypUTIBfRc38lysnKtUVJBZoEGxG313Pn3fkVnqpRIz8pUcqeLl
Fiuv60t+IkMKSw3OoedyuDJ92eA6tQPZ6c7e+z5U/JU5jRCLQYLDi8bz3wBjKGILiVuMTC58H6go
19YyP42pkRAYwd3aY1ApA754w6sHMsoaaJb8RcsYAZFESqGq/a3i0Wjm9yI+lpaXPmc7QhBnYekR
RWI/EyMMmiN/CgOb1XX+eJsuJQhRxYd/y/GRsgdBp70Dt0VhS0L9Y8ZdTi9ClwbFuLeDLmR8kzp/
+suMS2H34a79wwA2XTK4CzobDV5LsQDNfCWFOsV/n8hY8n9c/+VpHt+FC84ubwcvivIOQ7Z2od+U
WtOoVMPbluNJTwtU3ae+mqTsNoPZQZpstdhym4pC6eYwKVNMWU1OFf5ikS5ZHVZi8MgB9gCrlufv
DKr6nLgv1ZVvPjUgs8pine5lhsnNZ9cIM+DbihaZPLgUHTQL+UbEX+Lx8utmgmYk9/e45out1IGT
ro9ozavsNUT8M8kTvP3PsrBGSDPcq5X/GxmJ+lKSQHMq0rVXfZlhaec1wneax48nCZHb5x0yS6g3
3DCwH30rGr2nRhnkAovShsL21XCRe5UdjfKMoM532TQYg/zq4okiY1mv7kJ+jwlCtE5UwQ7Ddb8F
plwGwxHPlmWHWO1I4KjY+YBb7quXJLa45iyin5PF0QmWR2pDN04Uipxu8C2dg8BuC2M1O2WZzU0p
DI1r5U9lFI8BEYAt6dz0l4PdNnN/qmEh/w/NeqHaPBaJeCFeZ837gT5b2SZ5p/EacrW/NcT10v9q
EF8OWHd+h97IymStk5OprxhMfAu5je4fkNaXs8BznPPn+ziiIv3CaXXgu9oCOOPXbQM+NsLad2yZ
OtxicZFGF5JSpWEhP+osSYB9IwIS7GRnFqdu8P0FZl1TKCTrpA8YUFVu5rW721rNCz7GQNjMcs/F
hYiTF+ecayruTiQbzrOc/nORbDnGD7xR61PLWjViCHYLRuxKni9MTyzhvnIJP80eOhZ3JsAJvs+h
O8gWNtUv85QZghGENtPW+ldjsxH0JpafIsrMgIEkGahs6jBHLBh55MS8N3ZteTLMenreTtcFFqvV
raccGOzWGM05dRf96VsFOlEEkAahdYyg3m1Jjt4oWoyI+yFXWWMEh01SGMp7X0Y7Vz8qlTkGmm9v
WXl9SirRFacT4GndFNou/N+xnolADpLFEUehZlD18ePYlEB/sAIGiOCpBzvDnCKEcC/qtHT3zgnu
Lkif/9GlSanvzAVRbBPbgzp0pXd70qYJRqxtJrA8Xof4h1bFPblkpedZcqi76BjfoNVdQBVD0Zuo
iHF+mBNmCzGXPhxZ3IWPDj7XY+XFNeCavKjAvgyNZ+iRqNc1QZYB2Aa5N3oRdWWNpFb4R/juOtXI
2OZ2oZ4rfsXmcvmU+6gDywQD9JC4ARcuSwHtC2tpd0MnQSs7UXgu+rrnHvsmtBSDeZGmk8b4PkRL
4fj/p5hr0RMKHWIGB5hBM6rQo59Wn02uSrmpGUxED+VbV6NaZ5D9YhHc26yVBOP+rDGfWFCfc1rr
+oi2m+yr7CuwShDyxhU7O9RXzAmoyH9lSTnwpxUyb/LNOqgFyU/oSanVRAGuqQlFYIKipaJ+hIwy
GvAO8tW6oUO5fhNF1i6damLRjNllcw6iYhlx0NIH1SYFHmqCy3dcwmbbcp+4Z5QlMftpvlcV1Kil
A/v2EyDI5GhIExOK1QYWWq/UwT0rCeDCEm68w80BylOT9lF7bcpw9PFh3poRXQfVLxaSF9NwVjiV
oMaJlyiqZcCWBCSiR39eOJj2+uJIoauKIEB6vlzUqwY7uDZ0xyPhtYywfN9Q4unnWTVwf18067jD
2tVP1w94D6/6NDptYbGrf0d5SjcbEN3Gfz6TdyszW2WH1Av0edvJf691r2jiYFH1iKpcFnIW6KBB
1jxPAa5DTFLqNfEWN3cyCRnMFxwt1FMAA7t4sLmusAu9lUtFwKWWcZmmxlritveFxQ/vtu7hK0Yv
G4XbGqdwmdK/35ilJ++cRwDeUGBTtqgtdjkGiZn7wqCvGxQfwwJV9DPLVZ1HiUBCtUaOJQVg1nOH
gIzBe/1b/Ms+j/OCvxOuCf4K9PUiTIZq28eqCi7AUzMi64zQWGaLGHbJoTplY0IzzGZYgVS8jssr
4hWjerGweJ6hciyK0MrriEb+jgmsjE5zoELzdjPE0EDt/nxR0ECslH+Zzdp44ZU2qeAeQAd/PdZp
y9mFeX8sUNBBqoHRKk07PFzBSvA06lq/mp+JeBJ1/Wrvn2/23yqSlJU/oAmRkyVKY0Gp3l6hUCs2
JIc5aGt4e/siYQhVvXw2Tjm6LboduVlJbY95PYjBywGJ5TsDxyjb3csuj4zv9w9UP6xq6Y5Reuwp
CCXd1c4+kPpXGXsb9CXyakVIjS5/cToQmYrr51u4wTInNLdnC2+w6JTX3YNKSh5nyPuHfCS3oLwb
m8sVNoHfhdtHFnppJtj4+CknW1RztuDqfu1FQLwEuHcuqJwX+DhZsEsCHQMQMqoJDoHl8ot369l9
Zl+dVtEK4SMy1VEH44BsWVusIMyLLSVSwwm/6LXaNZYMPSURGxDAXvAdyJnLNk9iKT7Oi5fCoU+X
mxzgBXW/Z49S/ytEaeHp20qpG/C+0zf8Wj9Rv9V0N4eXRJQjEY75JHu76H/j8ipEmTCcLxjeubP2
UHnznCtW8Hen3JtnluvZCSHhoHILwNCeA5grIXn68BrdfVM7H33e3pAx8yXEpnV8jXVguDmRr7TH
tLGd8o85E6GmOigG1v7KXhjOeQBlQFh5uMHTn3pjlVVUDfgVClisjIwHCJFWTp2FuF2k85f63ate
hG6o4oi9UiSvTsaQ5FbDfCRNRwzywUOUouZdna8lDsidEIe6FzJh46Zw8bv8FV+LUf/Fjrcd4r2+
jKTXA0wkurxh7eJx/oTdFm3v4YnwDvszmlANG56aA6NAjMUq4OlGcaO2zWvpEDTjrhCNKVSQfjwB
F3g+3s2EIdv51Z/0n2Kmh8GrY18sDc1V9r1TA9A/6PL75trDyvZChM0Ky0mYwLHp1+o7WvJa/bS7
g6GcCF6hvNbVJknqgjDSZZ+UxxTwaUmxHMIgb9XiFfUl2YjUdK4+mst1+ZOXrJ9ZMKcDfy8ehSy4
heX5jCv8ss6ornlJGfzbE2wKmv/CztuHXeyqiV9ceLTUBUsOm6H52jlaSDykYCCQkNJgZVIDPoWN
QjCs9qbRZec+eFMa5wjPmNSS+hYnVC9t49/qB1U6ABm21wGwjO0dhAAYI6t+hA1pKK9ofqvnEdsG
9bDfZJDo2Ex6hLw2wjRyy0UAtxH/ObtZYT6BK6IGdOTFfx2kBllFwrX1tiPpEJ+AOAmk4xPUiHoC
gEyCjdDnp5BoB2Jt/G9WCQzI4dzfm425iEN5QP0sDi40ffTCDrqJYo/Upg2J3PnaviXje/6OVZ4S
qgkiNhmzZBrFnoUWOezSC3cwbWroo/YSzEnEepYVjGFyhNhNNU0+RyWH9TMORNbAhg/LeDBwt5IB
y09VQAdq34u9dtPc749eeeF9+hEBr1ymVzww55To2+HCOtgK0HJtz13BZG8isQgCzlDC1Oo7/XGD
/xmZCi01IH95rfu/ye1TvPWzJTnPLUVzvc24OsEm7/BFPWPECIu57lrMTWfjetTUch9GrF7WVDW/
L0O3ky+WFaCWYq+q7KeHk+NGdxv7nw1JILVenUzS6NUhh8Bm8JyhgC8u9hSIa3dE+Wo9f8FmsmTX
Ad/mTcFT7jUBw7gx4Yoalo/GqEnL6VsYgAVUsrA+AMQL3shJt17zT3C0g/4CKZdQ1lR4+RCt0iRU
ncMdjHX8W2dOfD7cv9p4VXDFn+M5GJHxnkyj2lzhE09JkbY4RhuADcutLklP/RtqbwCb33GoHnhs
/aL4sYSp2QlFMlJa9CqW1b3p33QJICIgECqWMJz9iTiSFHo17KFvUL6i24oD36AIfRMApYFBM4tm
CUH7uLqOBSW0MLzMU2vj/b+nN6BWMNQ5vsj9P4b050DRGCoWZwtZX8vAbcFDDMpceJm6wTT1M3wr
CPpCS3YFAuBjUnwDbNpk6f6AR8O/+gjs0Na1dwLKBHtVdOq2n64e7NSD/aYAVGAvgoiEckFZJw1q
7IgUQ9FkeYOPuGlEN5y7VEmlbqPvnEUdazejlzORNSLJkeaH2sIYeui1MrNOsGgyXh4y+zqEOjIQ
iANNMvcisGplTQj45v4Se5LKTeJxe1APsEHxaiw4L92rzn/ZV3fpYcKVDPFm2w5JaebaqiflnKef
FTvBA3j1DR8/CRq/Bx6fyvB3BPtFCq6Z0ioofXiiKRaBOMDBhJxK+zhsLIPiJQXMVtz6gdnI5TvP
6/txABsHCBzqHPs95xB9W2RaSVMioI8PYipY6aLvZ5GiSO/lLwwzAc5NEmyvZPukSokXoSgS/CDT
E5LOZEKrVPLZebaGlynnpl5L8oGGpt9eq/GmotQC8P7Zg4helRvfpTBgCxO1eiMZzXOV5ppaQ1od
XCfptEm3Nx7CaLcqiuPTlJ0WifjFj3dSbRupgL8E6M3CrNBXq6vL6bzT88QuAn9sW0MgcaXscBKl
QZhR0thvvcMtOMPhpNlli0nskHXOV5FI2ZRbCRATlhl0Ey/Z124DGd0odxDtJhW6BQYEJoDPTx2F
uCEMqvs2mltXNxIhyNWdYLchIFlR4gdhLyQft9fOwO8fq3EdYGqLh/mDtcHh/xjWd20Rgl1qH/YH
7FVGQHl8cFMpFhmbF/VWGaLeti/h62b/YjwV8SAXnXp3XCBf53FlAAPU6qu848VOEMrRS+9JNJH5
YswOPXdTG2dqxXCjiYsEYswLA49gFJuu51CsoU8NLcfSnW9I9tebHnw/M0dfXzRXTtEe+KsN5x5e
tD0IjiEBlHp8KIFfkuWNoDYx3H4pST3SmEsgtMT8WgVAiI+x4cyGZCeKI1qRj12mzMWBM6DaTKSx
qpbOIcgJ/vxcaAcUNopsJgHVfcZ2Hk5Q3RzjbsN5HYHSrUEnaf5f9MtnwmGrE7b45WjUlmzeD2Pe
Yai5Zk4pibhrpWg+wG7sjW+pwtLPiDowE7iY5z+UW6rEn5pPq1b7Rc93134TlIdMqpWPTnqJSaOI
arXoqGdwDGQBrzn/tDR4wkYAHsxZqck6iEa3kbdNBKs2SqwfOV3DUqNOEyBS+8BjSBNREwMpPMAV
SwsrbQwuA3wzr226Aq6RTUhvjUotszBGg/WXCmYjKTHA9TPQ/W5+4ZMPKvrG1VYacCSJQYAJbE3H
8i2OkfGSjb7yTRWSupG2AyTwRikiHOzZ5+Mperb2Fc0CZjNSHKphWgAfa9jgPqtRHBZXpYEPnlFr
zFnV1oRYjofa+6Iysr8KsGanrqFBa8loPbPA+j3dVtZUoiMV3ZLu2CHgqgQRL2YrBfePbzR5yG7k
iyn12wVlTMQgKBfewzjx66jge1PlXRILyhGQ4xCVanEWJXB0U/bc844+eeqDLOaqcO7C1UixwVys
jpKW+nlGwE6iIUl0lVeZBXC1lilEBgR5HEBlMXKs2WMWMeevi6pgRjbzExi20CzgKs+x0HZ0CG8O
dlmv22lb8p9/WZDGZ49ae+sjZ+yPOkL1Nm97P5c4kVALlL3mMlGMjg4UVA8o1mGh26Xa52ZNRYnN
oV1dIQga+KA9nH/bhg3H1tL6zkZsg5WGjwARPBpaULoEkgutDnBeOCR3Re3SKiq6LCZpVQT8cueN
hSdivAm61sxu8krhCJHrvZ2QCZjLt55e+DcnlMFL92zd5rFnwLf77dUIfLjE8Vi3S2QLBDSJhXLi
vXKkD44PcQ3QSrUvfbUa7d+AhaolwuwKtKcjOuuLVLQ1dU1L7fLcyDSl4vfWRga82bdcW0BVS5he
cGBUMj7uwz2PGJ+W+2agd5LMCkVt01szcWgy1HFfOjdtVQjYqJ22Q9sRRHv2lzBVYqmMQnFu7v5e
XWHwPpmaLcU7frhAmsHWk3IdNa9gZ039L1EnzVVsKppA2TyKa6EwfcyoR9CYZADGJMfmVc5GK37M
8rRyMlHRfZKNzcro54Z1p/OEfYW+QniZkG40FX0Avs2HiMxe8hjNFkSi4nXR2j5R4nVvFzgax+u8
vqQQL8RelIsuUSYFfKArN0J5sgMUDFsT++UWyn62wVwIolK+qFAF870eb0i4++xh0JYgNZl3XOeb
VUhqateVWsal//zgSXWqd4YjSrasWM7s3dR/oP95INEZGObIzhVtfKPWeHkXN0BHtLlGls8vKRRX
O/fySCmVP9nTPfxnjxci0NFMyXvjfnLXCdLpSvzzn4MXKjK1/cXxUC4YY/QSq84X/gsKgCK9Ockz
67Bv9SGOCT4sEpWJx1ixCkkeeyxyDf5MGqnfOoyiYXuetmD9WnvDxcOHkXwn9Xg6oanMZyh826Gu
EAx7CnEZmCnbHoId0sHnJW8OuHy/nUVyujwe35EH6OJNrqvxfMZGHyP3x8ddkMoCIuYw9cDICaDU
aOhPnDJu3HJFpSvGH1sl1EeP6TaKNIzdlJ1pSRjs0uk1LRzfLepppSGdOuTGBRcBstpyaQnHqxQ6
gUegizP13acA4vGFlw4b+kTF7gP/M148bmq6j/4mm6kxqExM1zqxddxWFG6h+58GCTwDpIHpELfv
bv5ubnOZHtVyYpjIPG1Ke/ueeS4PtYScPxhiRSmfr0ed4q8BUoHRe10G7UM3kRI3pxlGJUqP8pO8
Vyd/lKcX3dcty6BcRas4/5HYYmSlB5b352gRjKpPuu44K/9Yn/yixeRnZfmguKDfaK1psv7Er0Sm
RyzKHYnHSGbRgdfEvV6ffE3V5S6etbsw9Ihqirs59/eEtlw3CqiTm7/tJNdgUEBMFRhrMlI53KQ6
UJ2B2Wmr6AHrgcTFIu/UB7/lFjJkD16+Xuo/eYbtdeOEvD+CnEVLFsDACdbjahzUv9Y7yh71XGg8
Sg2cxhiJQMX7p+7N+5p+W5uFc3Y9HM56wY+5153qw5kUP/Eb4A03yWEXOcFiiwYeuuwCoc6MLksM
bo/MBH5LotnA2Zr4gXRlIqLel6L7w3twUELEqaB1pU4QAbToegM85UV2lkgjmj8KS5TlhO2qMjSN
w8BIvnqUB+ykOwDgk4Txs1rOLnc9rPk+eLVM0EDEkyxz7SobVdcn0DDo0kEC08pxA8xmLjfqJeYc
XFamdG21/TL5B6r+KMQK8oNvJhQrm4bFBQkR5HvRtL8VM5Dm7Obc6vPhL0iaV2STlw30RSCkhcz9
Sxt0WIqrbbx3a5ejZb30FEr1JjQNPMV2s/AJMbUs6V5TqKJ3WT++9tj4VsQZqjoXV9AVx8JdTU//
uyHOp5eF2VUGFdWsQvEuzUHVHxHMZn9/4XPY/5767UgqXZp/K9v6mAYtKHU0NhRQK55BJ8qv9Z6s
npScvdGVcAIvncXns+Zd7lnlAAf+pg2Cw9/3xN+FCFeL0qJldUaF9iZVwNxAe65E2mYUh7NMIXCC
KfhAmUQoMH/hVdgAz8TasluhUxPEBCSsTMpohZ36nkewCV9ZuD5LjHDFIQ4wbvnAYDz2PxYuKt5d
ZPvvHfs3/KDjhMCMuzA3XSAO2jDhWufhpSyx8wzszTaBo2H4MK0Nvtx4aJr9X2u0dHh8x7r2yChf
cHEXLX1UPDt9PZ6thikiYWwEFByTT+fk/tjp6SEVXffhAga0QFSfGjf4EAxahl4LYU0MMDtNAiLc
0oxAcmI3vKOrxNFibwh1g8EtulXGHWuFZ+aAfvBzC74QfRGIRk0QoIMlg/CgF48sRdRu9NkDdhl+
kTfPQBxH+GOXqZDNXg4neF9uygLvYu60NDaMrai0mOdhhRJxVYabpAYcsvzfcmV6GuWVRHahO9LW
F1JOChq8zqyNuyWNgUTKtAdAxAMTKyh/pzg+sLdlxo2j5pzrH/adQSIN1tzIEbATY0m6BvNRUngw
jQXCKjVQP6EY2LSvmgntiletw+de72I/JlcSjwQyb1b+YWAPu8f4Ru70b2KkwbtMJUX3DzmhUQlP
1n/ABWrm5tu0tAhO78s8AX5JMibv+y94aRQa1DKHGD5WE7wZO/n5IsU15yPu37rdaRlxZ6KNQwbd
FKWzYidL7OPDHlRDIBS8XW6P+7xeSTCJCLuvcx/VKictT0glFiG6v9OTTDvTJjdYA5GU6cViDMQY
1GpPF+7q+yRt6vHWcY3r0OOxbtY2SJreXjiHor3PdZ6ZQ/i+vifNI1ceEOBT2NHQzyIZyd7Lkx36
Wgu3AVIylUbe4FQitTED25dXJ7QabnYv9quI+xRKkBUUcULST+XBZv9K1cH5kJA9dLFzLhl9qGvc
HWcx2vToCh/1Hd0r6KFbHhDfchM7fmS1qW/Tt9qdPszqPmTe2MxCkJGoF0UfWyEYlJ36VfTb9fnG
+emxQTcqiVSkRi9J0FMfm7TqyR0QHJDe7s2BGf5CTNSbWF1i6yoBLXJbZCAyPd2aQK39QYSZWNX6
iEvE6WONcjflC1gxPI6am1CkYCOvELWhMUwwxGxIKuTZfVwdtVTW+RELDzIphnIONZqJHxdZswcZ
m5u5a3BZLcBXKXlzXoXM8Z13+5LatjNrv0LZf0TUA3cVBM2+BHeGC1Gi0kvrcVJmSlhVWN80gOGX
Wzdv24fa/7vlbjRkuAJYkRZ3+KonGapJnidJa0gMS3AaQB/who00YshvsDqlMrHx9NUoN2B8Nqas
6WDgsD3Kc1oKZetsRtsnElG7vFiuHucddbwupqPdrXOUuxT4Zjf7oZWOgM953WMiojUnj1DMPQdR
7bxunK3EwmwmdGTMQf4lTCUeBblx51u71z2KvfnV0ZE+ZH6rpB762vMubHA50dlOUxUQ3iNjiqJO
GhwtMXnJaiFUorZ5r4sY52TkeK6Izfp2FKhk5nvO2jjTimTxrCxgs5OAFYn8oq+0Fu/Giic6uuOQ
SZw51aQaugKF77UEv8FmqqnZv95imIjtY8LaGIL7yTHZhbuv0q0MTeRwa/+HzEd8YXVSwDaaS5MG
7ERwRGPpKMWPlvh9uRV+iIDV4IX9QEQNJmENcD/CiK443W9rLND545+Ppl/0RZcrOVhpVRfLjSlH
TXDS+WeH/iDabQEMkmBZJbtlx5VF9uIY3hTmlPqSTX3QDK80kjkgW6a7ahR4kBnVNOPJPxNB/gMf
MrJK8H5ajZIdzbJ4PKZhheh9qzAEoEGrvBATDM9Au1oYGAx4nPdMW9T8W/2FB+ETe7Y/wQhesBmw
vrmHHIbWJ1jjf2Ca7Lh70syPnJECwmV8tWGyaH8wAzzt7XTBT3dadyNjQq3/GFX5jcteUfNu+Un3
y9mqmJ4XUrnfwJEkzoO9sM5lpON9Zm724v7oUdtkeBviY1MH4Zkp5ySE4qer9q91Enus8pInWS5I
uZdBSmg9MJsUVpWDcWKsncuFUqDn7oeEhFZ2a9OG23aqT7wFUHZYFGBXC2LXlz9+0zszobA7kCZZ
7xeqPQ4r7eArE7b/2YU1foo5u7ahxl3iBbBDf4eU0eCHWRp6Y2UdKftmB/AO87vF3oxU19DV6rpG
Vz8W5qoop0ySFrIcvR2zi1yVvTa6rQKAVuqBSjt2v3vM3ypk6Fk5PYBZUH4byWjP0PxHxM6Yx3xY
5tuq8cjaWreMnpMtGr6AxrjYy5iBC8Iz6x05y+TTpIvqZwRDdDSudbsWK6Zny7oVkrnB1oNnqpRa
CeTLkIzK9ItwJSibKVJZvVFlQz7NGhcb9UzjGlhi/hD+3zj69om6L42rwYm9oM+2nI8w8ocWoqlp
d38wVatUUQ2qg2E5bpy5p3yb0F7A9wUWlNgB/XUj9stI/T68TN9nATtiDQ4AwQd4v25MbcBHWApQ
93SldK/LKKCkQTGyaL3qDWfkozB1HHPpnFFoyHSflFIBrFI9R9kOPNDo5T1n7QH071dFaWwpRxk8
xofHHv9Y9w+qV6edUk1o6oZI1Bbz/tzSmdMB4s3+zxtsT7rjceiXJtHDk7nmSMSxxQwPXYD8q5jI
jqaWd8rnhnSI0TASH31ePY8RlAp1OlUFLkTbpMGHAuM6OXwKhe97zlRIiq2CesanTaDLRx+Ujlve
ALQySb9jmcxFiTWI4L1TU9kooDLW7bPHbRK8sS0zTmjtMysKMyyCAwTgRIIrYGvTBOOufhXeySAZ
6PCQDA7UrjZtw8Qb9JuMXhQF5ehBVL7F3pK5G7Yy9UMGpHwbcvaDoy+k3sTrP7ZG+zhDxh3WLXhy
YkB+eaBiUP4+Exw8qzn5Mlx6FQeku7eO1gy+lDJuIKk8mauYEjKXEg9wAbe5ecqyIbSjZoh/S3hb
aMZdBwbuxUMS5BeMvxAURF7aInV43+qWlAqjtkhnXFXwcFtmoqfhvc3q0cfqsV/Hjk2tYpOFSOZf
HjNNWkmhTRXwxT6uKE5egPXmls5DJOp7m9OT/mNNMCshSzfG1c3zoc3isYPTPEb8v5+LyXPhNWFg
vqN7DBxl5KXitlX9fROlv3CHCNIF6YTxuRVxrk8H7wL4xOGHHBFn9is1lTeDg9PkGGVLQ9+9LvYJ
vZyb6p/L0ah9FngGLhPyReCI0dOl589lRvKfPZKzuzXpuUVQhyLpB6h5q2tg1i2bHarjAsX7eTIW
5hOEphzLD4EBsTk1Xz22K55YYGEAYTAtUaHvq0oOYxzr95zjmBI5PzKZp3Re6f1y3VIrtvyH6/9K
1y/XYgt0FfNlaoSPPMJVK8Yk/8ECYLUXmpRtuPWOxKFZ0ZL+aBFfGY7cxWeGPGZRaKzko8+jPwoi
fvzBVEpuKB4VhWiCcjghhBo+8PocXvZUCSHKMZEZtYZwGm9wWZHU+iEKZhIFS2eAu5YJtDBAOiBi
ctesRDDQJ9/svOJexyGeaA4QVfbN6cevoBZ7ykFErUWi7JuNhxq2JkBhEHbr5F5NRF4FQcjt6NOl
IdkUu2GT5pwCoI5i35KN+RLhYyk0wjxMD+lIHTm6JfdGuG6PsP8CoRB8L3A5+tmjKeSBoCFL3dOj
HITvOJNpb426jFUupYjC++3sFri081++wOHKSk1i29peap2568bOvBtH1IT5nQXtxoP/Dn6K/xGq
JLQT32CemRMYINUmjaXIdRZTsX8FL+T9TWXK6ccqBQO8SNkyYYmRZVd9jklDUcjP6BtronpMRgu0
yh3lgqmU6G1ykZqig/n+EXC1eCaBf5e0meftatVvkDQVVm6lqHkWbZOf1raXPniehSFrH+E8Gtrr
5D9SRR+U1PEDJWRBAR9aLm7ftxcQxSXp672F4TYNh1cWyBIE/iEg3VXndpqeUjupi0rhWGg3HP5j
5Lv+DkPDbkNh0DQxodbPDn13xLt97tupM61RjP8bMKi3pyycqHI+FYoiJgw1A+Z3nLK41wg9dGF7
yGBgqpNjTtQ00Vb0E3ogG3GFRyDI+KImOwCF8YcrgsJEjRV0xRNbQgG20ME7mXCloyZP7+OV9DJ/
knWbdQzQ51APSHWqQhyqBPex/raTFoi/0IyTLC0KmhgpZaesGN2UBfIpFH0uWayTPQ/wKT1cNo53
0kcfgu7rOsqtfsbY+xAWvWB/qXw/xug4GxlymKZE+dmRzfpU4pvo0OteXPAUWf08drOMLLIGePy9
o6uuotWcootkQ8tAwVva30CJEHRC9peYvm+6Go2h84P/Zf55MI1Qz7pSP/TPOgQxEk1Uwg5lKWIl
YQamJkZyJP0TFfKkEDRMNsW3M/Yte6vWALvLnLktyknCoiz+jLdEyPmaiUrf6K0UHl7v3y1MnYI/
jEsaDdckdInlXJkMG+O3nir8+SPPi9tMalJcUokgrHM6Iotemtt4b5w/4xSYBvu9ZypHcBLsNOru
TO+ZrRh5xDwMRjU8gLyjiP1yl334UKwPYEpq9J9r9zNdOUoustxd2Kh+cZfHdegckQtp9Gi0k+Zb
1baQpNimJHyceWHYgRgt9LLdGavMzWNKvT3hNsu44gGXyZIrwCKcf1nE9OxTiD41M0+X0SSATfsI
GNX0e9xtri9YnoooSULpJRJZqHEFCBNYvMEJqm1H3mMUx79ZoXZREm75QZXlbkhS6ECPqQ0uTd/U
O3jInyaqVZxgp5d7x0ECFGcbvAETRxxAgi/O8W0qavPsw18z43qnWxYiK9/akKbAvcLgMnfpQZE4
qQW1GrpqvtdUk++P4Hhiqe/oE6LpkKF5tYhG4ebLDfZg/qCQER0v+dHInsWJkYBi9F62b3behRVM
ZdHFxZjnOXBpwwsSmG6chTjuX4wTFHM48mrFGyL7xUmfklldY5peuLJ9C1wnxNZfe6w31EUQa8o8
FPvSwSW3pVVC8/S7xEzOSchlYx7BvOvXWMoxWoOcv2CjJF4LkVIfZowEtVMvzwzuJ+MYcqIrU7/Y
Kg9bpCcjnAz+1C9aajPXnNGkfBFK9aiiDn5RQtZjsZhnraRnwLutpX9rrNf/HM2yRinDHaswHdMq
A0JCWkikzkS0E8yLzaCZNUwiI6VAUAzaZcR8+8fz9SeQlqJb6v0W6YP+p3Os0EnIDwPkKZq2x61R
lW74qFWca96UGtGKuUe60BGsq1SOFwIfpp+MSR4CJi4Prd+WopuGcHXtU5esJ8S0s1oKJgVWvNMu
SIHTFrdlmWF6LIhdgHV0krg8xDz4JIWLC8QljqRlSj38NM8rH9nYOVz4OwNf8WFcWCdfaiZPtJU4
OOvyQ5Pmyri9zuc8fKkCFQw5B8Dnrr2oy4YDzoNEAk4JZjuPCNTweFDSCM72OqvEPbnJ890ChPoS
LI3Mg4gNzyTNVaRuwIY8lh34ZnbJ5zsrvWvYaqoJoDXGmJAGFLrVl+d1hsUbVbvxU3YpI7pLvBL5
rtGIf4wdulQdZvityMgeJpTB1cyV7GfHbZwJtpZ7S1tqvohvw/fhqSSh7f5iSlo4mMeAL8/AZcO4
BNHRWdD9TWKe3Mc3ieK0qTIa5+EqJ1uSQqnfWviknemMqpIi2S7ShXYFFFF/4COR6h2ZLFZ3kvz0
6+rbuNpApe3BCCe5EYfjrgmXOzoTuB/iWFfFBfxo9B/BHOYrYejs1qW+RJz8oxzX63srqem/ybYB
FXQTmhryt3IwjeWHrH6/U0G/a6KS75datcS9xvwFooq3Y85LD0H0mg2YCBQLeley13DO+d4vN3TN
JsS9iDMOOQacQW3nyV8u1Vz1JoYob+2UJiHyCWIO0NJ6BYOBtNItYuejnpSgxcyBHg2OIQyKpwMY
fVlfXeCwllR9eXSnxpFfFgipWU5MOX4tVpYtnZhcRQJPCUu4UKAPuQSMECDFNDl0dmruThOdJZIK
aaZkZdP3zYUWFUXVbBqT9iM3w5taap6+E+I+8EMxjEV7POE8PxJqcuiPCj/dJPLf12MVpuWIPSY7
9PJvFx8lkSCq7tiw18+YZt0gwZXJ/VNtztrZURFtxSrTz1ZTKiJ/3u35NBHIwOCcb1xCA3nXROMY
rQRwSzPlTZYu7gsOpPczhJ+Q3SP/hu+Jo5N06Fp01IvsgqJ+XRXVSSPb6L5twdVste/jARR8vAGi
/IlLL2T3s6p8uqL2ERfsKbfIc6tl20UvIQlTFSKRTrNUynvN8lqxPo9W7XpSx/Ri4o29FtA6K5s4
m6rYWlMMrcf9bRCOUFGv+TK6pqX3y33xfc5PC+KZWTNVMG7IyQFUOO+rsPiu6LSiCfRaquSkIV1c
zm0iZgaeoxrnDSSJoLMadeg1KWCZX7Xac3aYIHGXTE5HIw+hRVgTfb24BV+oqzjQ/hVn1v7t99Gn
tFfONrpaMoU83rcJMUeVwdq58Lc5OVIK4DjdGsRoHTU0A6TUi7BkT8A3HejvJKETqI3v9ulBaV0F
rsiePZWQypREr5nZSsuojBz/JTcuVaU2dFz2b6MBYvZt8qOVsN3z7AjTY80zH3Mkl9v18gPGEhMb
dfwEYEQuuIaGuITg6DXhgF3BW1xl0qtjfdw6DR+Yl765PMwHmMikVVEg9B4WjRE50wOata3ZyesN
YGaGJqhbv098EcCDUZEUew1ygrYmeKpxtLl7xykaDQYSevFKx9FE95WM8kmC8dN8RehA9n4blZWP
HUyYyDyL8S1mnF57OjErZ+wnW8t3mWNPwjk6ojCnFgBB3MnyoO+Gcc0XZvCUKUI8eQ6mDW3dqHDw
YBBwny1ypSihQmfwhsAqXDiex7sS4FnW81AlWsdp+5LjfLSjovaC1aF3U11Re0tSyoqcbFbIJ/0i
NEyH0eTce15/Apy8febBqJMKVNokxayOr2cnbyzo8wBFJdERQA6X0Oft+14JKDZ2OztO7GPNBTEu
ycrzQ5mIMyr/2A9dgK1Lq1bCPQPyPxghasWC9ndhaHDIxOcete0a2zzopHHEgqnJNAUJ3wwn1pqq
Q6fHfPHS31fQ+tXzK/pSoQQjXuSVrJC5aWYll9Pig8gSu/b8+4nHq0oZzh7RCnVwzqXBbg0rFZzC
Bt6TuQmIE8mAk+0/8STj2MhUiqzO/lLVlnm4KTE1WdPLqRyx7IJ9X6zyl4qWi6XcAnv+MgD7dNZU
qkPrJA7YOv/eBOKBBU6FsAB28NM4AYI7T8+w6k7+ZGGP8VvxXcx9k+wg7e6RbSsyL14UPUPow4je
wh/V74JPgzJuuiRXPHQVn/6BotHipDv72MuGVMVD35EoSG5CWBxo51ZV6F1/dAhR53eJ5DpPdehl
/s4dSi87+/EZyXYvxxYl2pFl2BNJorhHtnvhuTBk8hpxjlObZQn8BYjEOelZUBY4QfSzxYR6cssI
mWRYAkBoL1BZ9KlV3cfZOzTQ2ORg9iq1vFRIBY5xtrnAhpSMlqbN8zwSqTUvFKGF5TVDQ2+gMtNX
dShdoHO9TAzUUvK1Etsjy5Njosi7WRJab2PqZV4Fw05k7s8Q4SV7BwaIImUjjNejMYblcR7+y7+k
b1M4fi+o7nM9Peye5mS658BeR92Rz+kjwcIA9q8yFxQBZ78SkQ44wUB1KIqAR1yYwVwVnAF+IC3F
Q23B3MErw2dtpJJGsbb0h+Cd+4+Nl8S3perZ6TVPrqYAaI9ufZ6BigDtxyRblf7YCowGiWikFHfu
gLfDgRtygbZayFLfZJToXuKhs/3tY9GCVyUVKt1/Jl/8uRrHk7ksCCBRbvTnKDk9AX8fh2wGXXrs
vtmom+H9jYeFdpS1pTU8YIz6TKfVKN/yYEDp2Z9M729GFOlEp0eqwqoJcVQksTi1KmJVBROfvFyt
g4X60Itlb/1GaKoykKKb74NI04WHrlDC7khphQxJvhwZUtj14gRlYcbgfMNW1rF6TmfepeZIQPDR
C6NPwteiwyCVk4CqcK3o/vNAa5DSOIfzS77WtacgwmCnNTDtxx14pkbvhwjNOl1sf2XYzAoYpzwi
ANfUXKZwST3kwq6Y728GttHzwvGc2t3gwbwnzOq2aLGT/BDwyDbrBsBJs5ukbd4mc06XohLimxRj
UMByrAXrRBeFuBPnHsdV0xUGdtC5ejHTKnGbQP4u8NlekURcqtBrWlFfeuzlS1ILmUbehu1NXc2V
auxAET9o5hIbAinL3NrSFPQyfTLFpCgZOuFPpjwdZnX3eOEpIzTYZiVGlWfR5nP81gl/lXWhxzvk
uX0Cyod/YHS2fScTiyWz2N0E0hAm+6g9047oMZJq4Hi4zH/AyJtIeibzH5/DRh2oqGZIy60SgGvf
F4Q31xnZQJ1h2H9qDSFSSU2Rq1xC0373u/5TRS6bjlnT1WkZQtBvp44QvFHLZ51+UdNwh0zo/bVY
TjDasXqOIORDiokoaMKCPDjxCuiwGLKpZ6wgySGi9hI2PT+Z/HH1aaQhjwBSUfsNG0SBkfA1PoHO
JeX5JwC5mbdSeGqx+QOPKH7KQ5Xvjnhha+bJSUEHN5QxIXK+sqmZ6pp8jc73NQtWQ6PfGWV8SwgQ
5Eut9NbQbaAEwCAKlseLsMI5pSDpvIUvXYu0gVJBblTUOxipjAg1mepqpRFzE8HCvOAazx2LGBeL
4vQCzsqtv42KwmQAoOgJ9JSfw6kL5sJ31EfYG/zXeb1/TJAVta696HryHHsYsOhqKBKOQVYOjZUD
FxO5XXQaC2y/7szz5ruZyqPzQ/vAOLf8Xiwflp65vOrc8UDjP1SQrRaTpxOuikP9nwQMm8sBici7
au4HVFtK1AsBnrQ3xkqO2Rxp2fo12VgQJOHaXfXagCNFY22ZOIOnuvwwnpfTT3cKHLOWFultY8ni
+CPvsK1yymWLH6kGS4U7Ntzi4qc7FPWUBVtMQ5lIMx5X1mLZirqOF0+KaopUXPyTwhCddljuVQM0
IRwSr79fZpWpDxflLcSUZbzUJbVzvxu4S7kIR9r36fRoMIUWSZJjjSAUPJi1Jy4Pa+hmQawhzY5G
HbbNS6d/FLLFJx57aqnVqpu8jdKONZB1Yg4zquftiJKEbL58JbSHhGy++TSDWE6vHnuiJZMiyr2m
1ZIlUEoFPWu+LACvnFfqvem9iLo4htYTUoSFugAgmxTtqCn0cUdzzI9+pvnHZd/5N0dPB16d/0fg
8lGbwQ1QjR8H/RJuBHF1Px5kjd+gl+XXnoUgR6eCuB9F3gtmY+bzKWVd8auYiFMO1A9kl3SUm7F+
ACdGAB/mqRKhX1/SBeOTMu72t1taGVHhvGiTz5DsSIVjLF1TV0KGb2ruRCJbVzONNAn7suIB+hSO
4CYGVBc36TucEDe2qHYESPAmX3KWCBiCdTwY9pUP3EwBwmdf8/ybUX31LX/IDALjxznX8D7+LXpc
Uffi6T0pSc5X0+yXgD7EVTVHxgDpU4FaQ0vWq3Mxx0WmKHRIH+bauBDKlgSNN+DPP8PvTOvyHDem
BLG0QJA2r8SUMRFNT2d6IwiXIqIGA3ADzPvUBOiB0KTPTBH6KIofhxWdvbiUwXNpOZKXBbrwcM3/
nqft1AFIQm+iodXkRLA9UP7v+/hp9OTxKq4kzjERODGvHlqbdvrstTzKDX4b0ZRRse4xzpiIb9he
TrVf27Sll2KLnS9i8089x4jU4JGd0Zre3BQ0Y6ru+mx011Xw7WrvwtpgOpcpqWn0THLc/c6t1otj
Asunh1kh6jKbRZuW+LLMvscI5kxsmGEWgJ5iUpxm3PJNR+g1s7BMZokTZVp9RZBLwIkMgU51crWh
K5yYV7Dve0VSqrRqD4GQkcR9yM1uLcwInZUo8XWDIR7Td117F3ixngfnwug+QMsVGFnO5aeZT/Hf
Z24jJrJd1pCs5jSzeXiveOGaXD/W8wThiZ9o9jHclcM5/tLFvYojn/aP/TsJkfDeki04p2eLvKl6
eWUO9aH6tDjdSocERmnRDf/KoctHc7JCv4j4zEBo0vhmQCQ5iLgAj3wI4eg5IVd1HVaLInibangh
hIFPdVmxW/RNl9x73O78rLZW0QFkVbs0cy4NKCOozd9X0izp8sTaRYO9XwJM3fne+cMFlT/q3nD1
fQPKCMulg2b5oH9VjTRPkgdUXgT6u+fFjbJrL3cFEQtsUAYR6IDxcV9upsFX05ikr33DRhsnSfSD
BH3hA9krINUTBjRfsu0hGbfLZqtG1mCeTcGCwztUp84pPCe2ALYd8PzgQAegb2sHsyICb0bBkzrz
OSCIycuUtvbVdF4GYJGQrpSVDcwl029r/EukrAOCO3LWhkk/rkeYMyzKi+xtlEya35oJ1hx9OBB7
LzVk5V7E0sn8XkG/K04uJr7hmotoVP8sLikiN+LqkS9ZO3AqGqHzrtuGp3bSmlmPyf0RXskpkzAm
dYPJyFcBBJ4qmjqwDvkiW/2PzBn/TuhByz2OUg+UUPoRNvkNSs1PjKfviRG4ua8eh/Rdaym+SMN9
cQbs80/ZwtMIb5NLOfHflOza3ZmH3vk1qGJWpoZ9TZBhKEWrpSTsER8HEzJwULoYVEZ118AKOAp0
zhWFqtmvIRKewIp4C7rJWhP4gyFxIVGW1za/QUm6enZXuk49QLGj0neQMeV4lTsYcMfMaFVmzyPR
s+2lzDnVr7Mv0Ovpp7VCp3Yplk1U+p4VpNJ6LC6IqTyAEG4IRiwpK/los+pwTHzwUitUNn4ajdBr
Wx5144DbY8e49AT3eBriv+jgCnTIjC/aXpP1pxlg/3ZZvkadh/M//cGsF39NQTjoG0wVBHDDt/76
hI6FLX3igCVSDB2DidyJ7MzNWqkTodD0kS6EPjXQtbMYyqQ4c89PpThXnkOwRPPzADK1JqoSN49P
ztNwC4x4zJkE8HR/tnzCKjNlgdAfGUl0Hoy0ur2HBRcp2pZkN4ZwouNeQYwhXtrcM0j29qtHKIY/
fYxqC3wymo9HLsF3kbLGiDHxseYI5kHpA1ab6fJ6ElliiaS1/WxHUUdQbMrsR77Yvg9lwfFM0t17
8d9/MPhOuJtmgVaK1JuFWOME6G1FkOuvtxrCMTQ2/7Se6nA9kIwOFqnbjYUkjr/CYkEXpbmzXjve
Z6p1aTyspo8okIkUxTzHqJA9eOv4sZjLm9eRg8KRipH53wzazzAcaP8w+a9Jyj3pxrCRiy/hbC/h
FwlwoeINABei5v5MuWMWCvGIYO0X8kJOb4Eqeld2h5uOqXnffsX8BMQyLcqCaRBbnAdvzkO7GdoF
K+BQk3TI4Ry8kFL/Iqq2rxiNea5Ne0xJJ1o95iv4194JeHK6NnrrUp/r40yCP8IDoyHxPs5qnYpA
CuAK2doDU9sWloakbWehOZpGcqdiGCyUsjbUBkMANo0JtuxzYNeRju5Ch7qicZnQOW2g0eLblXZM
YqEpP1ebTFDemfl9YFfG1e+XsNughymt6RpFoAW4sSAQd1WJEWsrV0JKcH1sU8JTes5QylSxNLdN
BIMHx3IOOzuUChBdpNMXhyrvsP5FiZbf72SBhUsQ4SlH3YkNkcowmXkrZynlGPb6YZvPLb+GHcoi
fbEMM9iL6CNZngl3zVydHKCXZqqkH8IqzBn1cimI2L/z/hb1a1L9sVYyxXbQkQAz2C4YdIw2MTpb
UVk/P3dYBX/a2Gd7IysCnZEWyL9ywZt1d2XKr3O5LR+yjwM6vTkS2TvLlsD1KigOtF+ab3h72hA9
Sq2/YzT5DNnkSUvGaMXuiRjQgdDY8n/uQXSyzgAr8u/CayrgvrzzHbh2jHIZYE3i8Fh5iD8FJFJO
uBN8JFoZh6NxaO7e7TQTl0wGJWYMLTs+3FAukpwc9VlBDCiSaT1RaYNO0MZE4w825065rTMkT/zn
qLc30SkhieVglnx0q4RgfGMoKd81gqBYjcCyE8TbTUtYBXal9buSAZJ4Ysnc559wiT6TgbuZeT2D
ACyOyhKLT3ibiThqqM3cfcFXzEPIFaIn8lX9AyVTSYVYYOQRwiRngI+K6tKz6GAKNMJnL5iuG8nX
Vsr1IH9PFfW6e9/Dox5epiiJMkSQKENNWHZq7xjcNckHyaQOvlC6ONaV+PXJ2ujBMy4cxp8AjgYl
5jRtPum5tLSMQjFJDnpUmqX7Azlq4RyQqg4q+Vuoj4Ngh+I4ztEgdtBVSjFcmErofoDzv2ZmXzMc
fXTf5+o/GhNSdpu60q9kaF3MMw1/civ6AwQOU/2PuoDD1sA/vwAPnPoK9V2nCUifveuA2y0nz7I6
qQ45RBEQ5PTTQQqy2JUthzvhFnSgY7+pbJVLD42GbgR/9cUj3Fv2Lg4k9KOrtmHudV3ZOma6v0Bo
/y72CeT9ISjg8ClSzabM4EDubsq5EQwDDHH52CYHRJOodvZlZE1mlHrkLPDg2J/8cflg9ry3tYdY
x9F1zNTVbQcf8STdNHoDlHKEOJXcjb1Tap4K23SbAKoM7E8joACpCeE5r+I9Sddcmdc/GnHk7u2l
ZSR8l3uqrbE+bK6wARkoORGpHjKhTkj6fxDhdobHUwU2uRiCntyMraQ85jh1Z3k7GDy5903Azah1
1g3C3g3YZALtuHO2ODQl8WdYOhmyqp60X7sDTXfLf85Kszdpb+3jxH3SdVvBcLrx8VwufBmlJbD+
B+SElpoaxlSWt/mLW3ZSmOp3JKLtzhOTgwHxIalAdk2WuB6TcsITGk/kmW119d/aWN/a1F5wUWUg
lLAy/U2ZUwKYCvn1hFdr6bPDYacs+2/w9gebaYKrQf0TLYBTxbaPwejjCkJEZT7sKNtdMuY9n3Au
HT20iWT2V2rPDZxktASTb8Vv0435wMYSpg5AECujlNhUjwA2epd/LIoPKSiGEKqtP1Z2XhXHc+N6
2xTEF0xpK0oTtmkm6qQ9jaERwlu4NcZwerd7af/xj2fe8W06ACcuHaOYedfYqg7pS6tESm6vmhwD
jdozSHITY45m012zjt3tIfFQs7tDye757N7HHOS0r+5Hh3sSbhwNLoz/zFvnDigvt8Sr/WNdVP1O
Q8RcPXNnbOaYWDaby5wbkVDYb4TMJla7kTbeDzoQefSFyFgEIun4/RtDEM7H3T4mxFCfQaw9C6aO
NKqcbn2fSn3Nvj1KQ/bPNZvktv8MKL/GgupWYlO8li6Bl2K7HA+HgIcaR9S3THn3tMe6Z/OOITdv
KnSAYIWeHLyNY6LLRwLB+CnI0Y45VK5Ip6O+op1xP1ycFD7zkA9uhlGz4NQlbQ1SfmLoCVMBLtIx
+x+KQFXAja0zcsmcQn7SED7pxahQ2uHG2VOLlxhcp2LEwq0/g9tAW9mbAdw7WE4BIN1skwbygOFR
OAenou3ljM9rDbpidsJhA6EwcnjSw/6RYg+hjoUjPmmGO7kRNULnqOl+Wk/rdUZQMGAmj2Rq2Qum
MiA1QztN4KToLcKQR7+8v4gX37owk9N+4PmhKP3YnTKxPS9OBkdEN7sEPexVfa/w4uzOsJQxkY5l
SzlJT4Y4CKbBRIIupIcHD4JqO2lo7nEgk53vA0Ns/hzC8pN9E14ocHvCUCYnwRxw21VVBGstKjZx
Cy2L6GnpD0CY3qyHI+K2FEPgwMvJ92xeB08jSGg+8zcgnUBGvFXKRUkW1Zt+63+M1NyRIMstEiHS
fRSQnTeejyX28uGujhI0AmXzaKISXQZQCidR5WFy8MshnAXttXleKl0aDeir45LqyGLfd59Mo4NG
Dx+v/YqTd2rbgYwpsXlYDTfs2ZNuTTjIHT83+uBlyNEEF2MNlm92ey7K7s0Y2h1ZpP/GIeKKvsAo
2y8QuaaEL96BhxfghcFvQHeQwBUIoC+gPI1dWYDqutV48qFVRierDR5K14OdJQJtGtcKa1NoWqwj
RO22PSZnuREQJwy73G/+PbSmtKepMktWLSe5JC/rY2U4XqjFyZ6605I2TgswVSjJGcZZEXeyQ63z
cePJ3oFjU5QoQHoYmnsjgmZEPgpO0JvEmw+Lv+5HGXixk5v4Rvh/WWflR+cqcdKXL5JmTkygld5t
BRX/CxT2on7D1YM59DHCE+MCez9u2DOJwe7cW5rRXjDYJL/6mmsdZAFhbkDSFgfBTkfH7ZXFwuRd
m0Mw8hFtlUfmItI/sfy39xikbPJl+sJNEWnwLaf9qlnFQXtJ1LI+NEZcOyDwVT6x0iXsGDm3uATy
Jj4wGHEp9otYNd/zLC/NYN9jQEvYP1GV5bXTYmluruMnTJu4cEB4ZKsC+748Jal3U7a2YSry0IL9
BFgqIoYpqQOyx3n598tsS/U/84RyLY39xV3yGryYgeLOWdbQyEIDE1SLXVTCNfOEde54lVQwmBn5
07bOh0XliHsw/15jxoxRQ03lwVLFClavYqFFYSxpSr9J4pqBv1iY+nP7zOj+S3sEJGUvtAwPma4b
yVAprmL3FKz/ASDgHSMqXQpx0+uC2SMlAyDNbhVLNx3X599KiGebqbLcoP7dhQzdi4rLuyAbma6p
0jDwmyisHO18Qulu4wrlEVHl9bxRDID5n+hpoR6MbcjTy21oAlx0BGs/GAWfPyf0PW2l1zjHfarT
vlasdfVFUafRBn+EH3odOQh50IqtN2yWYDofACqUJGd5kbskuHkpTDIP4xjqRnMvHaAuL/8zV/ZQ
JRmQXm44K2xlN1FQdLcRSuqifxeKybqHShQ/UM9LsH3oQcjIhW3iLN2yAk6AobbxzfAJLg6gHDyF
pM93yLAL7gCAHHEyNC795MU/YNab11VawSabglUcGAKsFG7s+FBaD4OCz6700LuPyXsO+e8LFQB0
CXDofqPf6Rcw5CLoR9HSD+PB78QFi8I0V675hIivBS8EVyA7gioFMWu6Kgc4CMeAOgFpsm9aXZx+
THemp1w5Q5I85bGjPedatp0fkLzq+gw+lTDqDtojfRdQKHKy4BZZjl9V4hwL7RfADtsDU4PMBaH1
BGw6s/rjCmqAFIL2Kho2BMUo4GWrE1YCyz1x8kk4NRyU4Lu9mQyL/BzLUfUeIixuIosjGECtwbBa
hlB8Mi7NKrWfkC1DbuV7oE3nhHCX1LE2jYw/SoeVNk7C0XoHKUS2fIEqHUxS6mtaIuUv1+396Hzl
eRSUZ3thSdNlyKW8k9xTgq4pmcz17KEYpHJCxEdx8LR8p1EbW0fO5ePe1SSQzK4MdUtPfTEM99En
W5LT1iJpFUyrxMUwFYZzOu3MPbYGC6iqRqLAGoy0fjtI20gt13I54JnrAh69iWhi8yLoE6W0T3je
iomxjVXYgGG8VEXQc9qFfz7ydGIQO6XjoNtw1+cyGK9G84o77Oev8ah9WZYedXKRxPRVg6GKfu9Z
EiNoH4JL27C1cM5P+cH1AU3/V5AhQBV3dTt10bXitRyGBIhounlHTAsf3NbwNmua7/qh4dZR3tl4
LAR+M3lVXQD3/UZJA8A5AGiIHc/1rTifIvqcToIswDK+eTvM5urdtbh9U8H32hz9oIjzM6jIFuKV
zCAO/u209R2BZX1yE4DWiXaEtzpHuzRBYj2kr4hDepqrZ0a6fVkwyDDscyX9dfVpY4tSs7GEUZQe
miM32kSxwaeZQhCQ4qip/LwvY04u9wpmOMjvzORpSP6dosF/v+QfKjWEDpb72UbYUjvu012c4Mkh
tVvrTvqc40sO358YgEtJpmto7xgjZ35MU7q6KHAh3Nl7vmQxlHb1YAUkbInq8hfI1nba3uRxrHlQ
ItVVIwPT2er+9CBYRVD7Oo2Yw3oE3qvkcBL65ANS3p/qVRjlEkbc3DRMnWJHjVsboJ94LrK6VR4H
cfmbvjBvz18n2AbTfcelLq8xKCkfVPDiTdCiOF1ze6nD5T/baR3RNy0wwCGZaMRnBFbQWguq8BsP
NUAYeatEz+OGHlXtG7s4tRkxxavpJLoxvRHhhOTc9/oFKSyzEryKiLDvPGj+PMUc1LA7/NeItiQ0
nmlFVgMhRFBSmDngNtodQyXcOTUYS2uYSXtl4Lor+Or1A8l+1A5A7JR3YdDxGrSnhpV2WDwKgEjm
zFCZgKThOVgiWeesLjYlS0nyQoDwVt49noHRGhxad3PXz68mv6XK6Wf+juo+yt6gPV60bAflfXCt
Xs3jx9v7CoSdnsJ9x/yjAAG7DcHATFoSiOfA+Kg1TkNTu/nIadQJIfANSz978rMG9hoxT5+6PP6y
/pp6uS6FjD4scZ7robukect2uNoCd+WurIEwscTUNtNKutAtqPe6s8g+vLvPTLHV2AI784chSsSs
GQSdzm+gc4OlHewvwaKpRSMd92os9boLmuBF/l/x+Fy4aQ/+6o2M0yKkEZNO9cMUjFgWyN/1J8VR
Qv0oIkSKiuqmAQvYtxvO+MqIfxLU4MOrLbBTOG90fbMtTChJtUSKMEBcWooQ5kvRdrHcMHzuBJhU
v324xuDoSg1oq0FAXOsu42Ali95zRGx3T69FuQw2ut0cP7aZ21rMNyXZgpzxsiWBYxXp/+osBKB/
c2pRBYG4dXUQxgPyEup+wgC8Mfpj93+4iZQU2zanrf7gEdILnUMEj7PizRlkQOxl6fl/lrAGu26Z
vszAs0gWI+ye9vHjdj88U85NLvkqjvPWbRBSYLTwU8rS5FZDI1ovjFKz/ZvXiBcWEZnTdlFFQ4+A
wRbD5VFR/mFZhKPn9nBpD7+fQgED0Yr0ZNVe1ssrU7J5r9/e0Ak2xfGuMHP9paehaKKVoLDkxkmq
BeVm4I6fP+E8XA7apcHRiOj/pbbG2v01U6CETyZCcZMW/IvMpzl4gsrBLBMM47ZLl8i7+Yul6f7r
UK3VUadM8VoNHn4KeZXGElBRTzERlYnGy+T8WzkHH/S0uCh16Ju6r9aCip7fHO45nMNlwaOlWaAE
oxH+BqTCklBmuwKlv9ZqS31haRT8b0YmXzH3wn9Barj9cV7ysvrTb639mvzNLdgWdEZYruKyAto3
in5hK4j/kwtJs4o+zFOR21rM+qhb75Ovpv1LbYbxtcYRyP3pHZPNtqWaxJlzsNrwEd+EqA/YtN++
+aIARo0RStn3DAxmhIngxmvNv80m+zwozDjDyauS8/AqrS6kz/dwOwu6JI5oX1ux2zldiUukGbu/
eF0iuHwOsIXhCQA0rwBhkYBaM2tfibdNNH3p6zWnbnDnI1ZmbEV93NzWT0R5mA6CPu4IIchFZ0yg
M1SPQ0W4VvgDBhF6tWewrEJv6ApDFSE5MGPyfy61f/NR4gD4rzsmTT1hSoWFknlG6ZDEMmUMI2hv
3rZfzG2S+iHUyKhDiGfbU1hli4nBc0IU/QuE+I6NvsbjcLspiBUlvgZO+kYLcnQLnEkZvQ7Eas8B
y4hzf1n7hWuRnUs4wTgS9rISO0XtIVtDqcdv1lnErP7HP9JId4QWqhY8Cgq7IoC0Ymp9spkIynKv
ec7br7epBOlcazRd/HQeH3JSQBLsczjWmOg2iMKYjdjyytM0WVnjS5Q8Kc6453mNpqmGjBK7WGcN
sXKpnI3XC5g/Hy9kpEe9H65n7fF3gLWYSF0lnkyTrX0pufJwmCvSKrmsxBiUT1TCFXqSFgcQKCdl
78i3G3S9OMUYAYwHxnvRX2dJc9rKoxs7BOQbzSfVA4KfjfMvUKlU0zqwMMTU9AV6V+KvouaFIkY3
oXKCxLN4f8Hw/TqjSPk7pKXQNRUDPoc1A3EMRGL+l93z6+XDl3+IDF29wMCpZhHov+0U51u8AjaH
4dqqlCRhK6Rg0IRzAOvzV3/euI9lEcDsiwL5lTgUQvHNMpeoTWw79Hy+R5pVJCd1AJfiLifDgGqI
c4PkynI57atjeoNm4jWPfErLKGeAiAT7AUm7nSaPbUV2qZ3tO1d7aeMnjxdvMJbNxlwhQSiGZBvM
SOKccuhIX9LeP0DQEWh9ftQAypiJo/yZbUY50Vz1QEydM6hX2RlDm3oNlRrhGSAId5c4jQvA+rZe
Z/JucdsIpuxJ93ZSWnrS5N94g5dWYalAQMj65VwAxu0lE4b2FXwmVly4YZLZIpHO8vAMdkUCtpNz
WoeKWYDShJ1AWXkWkzTGSiku2nhb8/WTDBxZ4HG6nrAS3gkebs3dQMwB7KjIyGMAJU16G0UTDnES
VoMXxnItFKbZUuUi+zqJt8EGAOvLRKmZOVsCMzHsWMyQbNO4TFKRbdHziIMwnW3ycFfx9X0+XxnM
V95USd9qRov5hBw5zK4m5kJObDa2aDsdeQqA1xfYfqT4njMPqUXBUL8RrZXKr7NiPrgCf0b9U5YZ
TyaXIsjp3rxVAKDyHNFx6FxwEdkKVkpeFWEXh82xsuKoUePn87khGNrX4x2x2dFL8Nz1QIpsXlxm
U9mHPyPnUlS1wDh1CppiGbrN7mOgGJO3+fCjfPLbI1HxWglSWbzy5KiuPEB3fZau2qJpxOMJpJPr
GImJ1L0yhUuQa0rMwKGKr//89XU2PiMy6qIG+/VjnfCRQtv2B8K5Zj6/O44EcaMn7IcW+RJIVRVq
dofH1H0JzPu+4PVYo+ZoZrGq1K+6W6sSccUufzjq3g/4Wae+f9ZdwKHHPRYWX+ZwQpnT95x8pO76
Q8z0ifZkq/t6Q8+DlIqwC0CVuHVZTeKel5ML8nJCDsvK9zq7tefIRdGn+g4v7CEuqHRmi/HnV/UM
w/ycq2gtjmoK45HYK4Pc+M4p57pnoiTdZwgKw4G097Yiy9s1a3vQu88RU1gf2B8DdoYSfD0ZBVCS
52FzGfBcdAXHLlh5AVCkt4tANMpqb2A7m07iDnAj+tH6gglbbrPMTr+LddUSdRzaNQUMOH7/Zxro
btd7p2FSNIfrgNkFUUS+r6Vx6ET5S4Qr2+Ayyy2fKkp35CDLCLlDXvpgisWagBqADnv9bgWloWS1
rQjFImvwC8c3mKIeTILL3qOkoaTHeaeOqfXWmSN+f0fFYO1Zbrf1fNuN3Q+uwmfzLpP4HmjuK2fN
/87gEi8EiBEZD8ZXTvMNhKZYi/Rwz3NrXdfDefvUN4JuzNma0KDj92dYL5+aDsZy2AbdmfcN3qBE
OT+pC5uh3ZKOqb8u0PllcwFUPhq1vBU27Ew+QJQjnUYb+pS7X7h2VvXIue3H/9GrOnmqp2tSujaK
kIwCozxa4JhWrc45mxDydTkeAyX7UzK79q0wQNd2cNWKFzZfSpw2fVZL1Moso4cId7tB49L7A+kT
w9oXlqWlsrzWDcJ7DQb9VedIMjAsJzNV0lxEecLJZEHSrSMjP4KrYUTOrpks5Ew8DCfrSauv7H/0
Xm/agFmOkkPrVDX6fqs0HqC6/qHtRcvMxb0N1ObVEbgHW0s8vZSPk2oP+CaIahGDAK5mXpLNJlXY
Qq2mZcBUpIAvXP46BVJc0T3ZCrbvmHVT7e4ySFqQvZjs0UDSImtoN9NKpjFUGHjrZdt/yRG7UW6Z
XpkoypUAi48/uvCb4ycqjlHSNJ4IWp3MptwUgAO18wve/FD1S5/Aq/xsjLI9vXnGy3vPFBIuyKr/
mrnQu0oapU0NC/3vVlKE7XkeZ1ns3JmdlYVUXflAXlD33YhEF6EQOrAyzV6gxHt3pHy78tlzjtG9
F5ukzssDkZNZKSQV/KBGDDADX3ZfWBynqAA8+pYT4QTO0R7tyAEAifDqK1CUnKyJrRFCAXM2saJ8
Dla3vbP1yy2OSurSwgIWjEeoKpYU5xXguTq9Naon1KorO+9UziWaZ93NrXYYMzudDDTyljpDDWlG
af5XyPO6C1NEPeWGLQyCOIowfMwWW1XRJ1n4ZkPoL/Q/8fTKRc5hEwRdvLkWN+39vDRhyNEZDNmX
ewAk+H2avLVTp7QrFhhrgqazULZedFzkv3Twl3rRQAo2Hy1phRA9MVGhNbPmn9yQvVUlbU+Pc+hn
AMWJEWrI4eculnjRVwiBJKtJysS1btaaFo7sB6DhLdUwgRMcDwGsEj0mhrcNnSD7fM4gUc2bDtbs
OP3mqfanHN1risGeNMIVbV3jOfUBF41pzNMzN+lhrgzKxmZzTAfxJMWedombWNNk6Yv6Mdvd8VGi
2FYzyLXYhRi2XwewQcuYfuD32PUJCgsFAXkdqfSebaUmFNYw0SJ3MwRp0k7os3mgUPvdhsBS0bXz
RnigoF/vRTYFrzNu10dTMNaEWwtWZp7GHsuKW6kbVrM36UOI4wpJCrcIM75yvLRQ8n2d2z6uLC9M
8aL/XhFGTv3JTZDu1GnjN7johTVZcrwtYlFIhj4QWz7v13KkfUan0ZS0PUyqySLx52oB0P4c2DAP
HH6fuSNbZViUJyryuP8MZyOPzJN6bWPIEwhx83q/B3/kcnF1ZEZOIH+3ipKd/ae/9kZCh2LqhVXn
AOQGTQ5+SnC3Fo10kAsinp7jR+fEZSvZu74FuzOvEaGWdhq3m7Aoaur2H6B6uhO3oZwpmC47c9fv
U7hOLzMa8VNXNR9MmmdVl7WKk9WTtOmLTUFP2XHAszF3sAP1lYfOKPrb4YOn8kDVjEKytxOdVxJ+
ilcX2uPVNdgwXOPUDA1nOzc4QftPZXH+SFU1W9eceizlm5FtY31zcuGgSvuS0PKLSH5EGfKwBnDX
dbhDqaAmhhNSvDJ+0fmomm4kMbgzQ8LBfGwr7POSLYzjFgPo4JxA+DGf0EdBNjcJkxyp4RFAB5jT
rMC0gTiYv3FeBGq/n5CPZff2LgeiFLYPL7zxMCxZo9hTOEc2+knynGM68mKaNXqbZCN/YlucqZ8o
pv2z7gZlKwDyCB7ClW7H8ur+Rf+P+/qzI2PhMV8JAwNiomBiKfa6QRYjGgVbVJYC7rjsTXqbB3Fj
dngBdquJLpjzLJG2sk3xnmIcY3S77HYR/CUNpZt5QGDJZBV/x3HwsPm8vN2vmkmLkia01AlsYF+4
kkcU8wf7/hzeyk9a59hXgz4mxw6vP0Bp6tUKyQS3TZ9zhN1snLKw6KbyWkdipQNQYcA5f7kUSSS7
1RrkH4osAx9kHPHxOuATQur/SwRn3OMlNluHDx2t6Gk6p1kjRKaA8AyO2a7RPXISqgwNpiehZL1n
KTt8AMXWCT0iUS+ZsJtab63z5BOgb8uZwduVaKlf4Daec5dz/l5OzCieAX73/sFU701gaEv4diC+
V7235OvZptRq2UejCAbsCc6yyT4P1OyKn+0ZAOlHwrHa0zCjJmSJMxu6Us+tbqhO2nAh2zOPvaHi
a51Vo7xkhLgFHvXhyyfWlpW31jIVVQFh+G3Fewfc61Cck5JmddOB/BvU8IsO6iUoRWwGZI8nLZci
IRtpALqdvHArTM8LjmbSCGNDBRNmRRN4RlCKTI8L93Vimd8y3z2e8NGiF6w41PgC8oYzcT7YtSlA
QH4QQuZJhuddpwyk0utLwO/aNTwkPGJ8ZxBwY5uJuiD4RS9yhaD7wgWDVvfB1bXs132NKa8uB6+O
dHudSy/mWgBgpMdqkUuqQDcet+R+4+wSoTuXg0rFZ1E89yhVbcHRDBdVl1exDXtjX8erGAAzxgyf
blNF7TOTOWMCvB1whP8w1f8sD5EzbpMhSjE+11O1y1EIcaAjNJkLsBzFuiWyiQIM5FtEhYJmO5q8
NebiWJRyLdWu9uveiLkuSJwVVGb1wfr4igHAm4yyBZAaa7odmzcTRRYmxH7l5KZuExTGV84Lkh3M
WqxBPlAub5GbUaLK9dmqh/Xbp3TRQ/K2VC//NZeMnHhmXhoKskJambMF0oH6OCOqOMEdZo+MJkBO
MoHC9rAviYVogjmtk+nVFtlV+eKASsrBHqYEUoFP0sP72kHKj0sXPh6vPoLCZIu6I3q5OPAicVyU
9v04CHTY5HKm1Nufs9Yfbcalh8xIPUZeiiihrNDmn/vsSXCpL7COQlNUT8v1yH41+EsFWEkIQ9Bl
bYctcioiuNFD/Qvd+XAvgr0Pqr6dDPUllKclObPUZhdDxALkK9YQJsfPkM5O0ibZMlSsrqJJA/iw
d/QbTKmYIHdszVGUKH1YlUAqI8pShAZfvQfTgwmgmJNKnBNvabV/V5I85oe/u/av6P6skHz5SrKk
xNgEf5HHwddVGCW1EpPV5EXAafrwuwB//GyDE9oz/FDkv9w2UG7QsLHBlPR0od6XsyAMAC66oeJr
FjlZUV7WE2uFGEwMdMUSFu2ztYv49tMxBaEa58mCGy++UzJaGn78bBaqfPWmROXwUi3VUSzmAVNm
86W3Ri72OyP+hBgI/zCHVpOwVDiW/vpeVwGf6YP9rMg+VXuVOKLo1JqvaPS+dtx3cZ1SNYo2BZsf
DDAzjiFqQVmT5CU4l9cDpvw1E/+oCifmM+qoiiBXa82ODMSAQeLHBTFyJBQVHKL+V0E+wA+owy1h
eHv7k5Rbrz8Yxs2pFwyM/cHF1IZgb/ruTuaD3z88v0ee7/1zAoloMRdeR+GbEah7iDzyl5Nz+3Rw
LUt4Dxiulee8lQVsdCoM6wtezdQz1zPH3u+TaoyjMQRyClSy/RCJOQ2msdjUB98BJMZeuWueYDlC
t4/2sbOVsounWO4EFTr/pqU3gmfa3njb8PFeZ6UUpe4f5XoFF2Ah4Sw59KTR5GT9JjACNvHpziax
pILCmDPYHonUa4VxnuvpwFXWIRQoJXu+6Ob1/AMxTeNjxM5bWPT8yH4ZbOfVp7TRIQ8MvFYIoVLe
roPjyshvMWX2OO7HIuvHACPOuV6F4VMzeLlsCvNtgEwS3OlIl5MVMTojRKnm4SegYI5rvo9SyKao
9LIt6mIh0o+tNky1mcQlTpbKREjVj44x30MKL+ArjoTPWaYK2HPKLVAk57deyz8qSA2t0e1S2q8A
BCDTUh3ATpi00ZzWNEO4rAbrDbBBQxzZFOy8mXXMOKJIfMuJgzWyjYNTAWR0dmLg4vXpu+iUtQ3Y
RPTuPFEAenR6x2U+TphL1I0Cy5h9/p2Zk+yywkgJiWqT1MOJUxfogqTp12P3sG0EBy9cAym/Cv1a
lqFM4l0YLlq2x/8CqdxVAUPfO/NWS0s+yBhdkit773XRoPCKSlbtx7JNT9aIhpoTnk3vuM1L2wbu
wW/ngul2Z9vWV2gYRsBh4SO51/PgVmqAB1uA/9VOpNYlI1/ptq3NbiR46T6C9xb6A2Ttn0VkCXdd
OcoSBli5GvHlEhWc4iiJyrG7Yc9FmRBNPyhL1OOj5YCouIB4A9CBR+IDTZ3vTSizLpilONfdrIzv
BFZHsWpZzqXN1boKbsRdnpYPIApSyxuj1ZocmBG2DualjvWrD5u402n911GjdHN5FRVObBhsikOn
yr17ge0qo1JofZn/s9/876mVceKRkfm9uDHEGB/NhOGHM5EMTM4Cwz+918q6tGuSDPnBVpp2HXLR
koT2GA4xMDsrOy+BGfYQcg9kgR/c+2cLeKMe1ujeMYboROHbn1uKGMI1KGyOjUKhHOLFtBcJzhwo
JdKW195aTiz0A19vPbPM7rgiJ+4jcnRp+PE4AVnZyQIhP8HsXTBvH4eukE/X4PNrulOllkW0lPGa
cJQoPn5UWFSBhGAnr7lGq1UbV8LhNP6KePrfzF0SCbjVPV4lNXWxdKpHdDobylw1zOfKY3jWz+NW
dOh+asosq9F7lOPr1JFEUSYTCUrjGHvH/6DPHDaqKND/LRD0plrPyLSTh0Wn4Kl+KsVttn/VXnew
MR9XysEnK/gG4QrYy0n6Yg+fMjXR7ZoxgdK9fJWKSpXZG0VMxW44y3vdi+yqZT+/KxRhsfEk2hay
LXK7HAXcStWecWfgUqtq6D02OZ1TiWIdQg9R7p0w0Kzlx1UlPrK34QolZin8EgdTlgETJ4Eoo6UZ
YTm1odMb4qrMCRFqyAPLyPyxoK/deBvq3uSWVWT5aqV9Veyy+ZbJSmjJCyPZnVdMBn3ve/4h94SW
7ySWzp/VRJkXkOTmCkBBDvXXvdoXK5liQDllqoJgMOhYs0sIb2kdbJUDBBI/81rOf1JZIt74m8ML
0qimgF1SzAKx+TiMqU7mRW+h3k5Ads/DNO5kd1IbFUFOGlJWcEoNLksZxyf/JFzCF1/1HpmxxnwJ
EOwdj/6lwlEnqt6EQMKuQ7sAXkWi8Eq10KQZBJlu4NogFSuC+y23fa7zgpyw+/TMQx26JQNn739w
F+w08Zwj4UHFo514juv0bs+cWWkwZ0RFMtAidlmbm4/dKhGKhe1dSHRaHSmFWTIgSqZzmFIQvKAK
s+fNbQgBKSfoFLYh7gEZwtCG8q5IHARE2W16d7qJvZ/NNvq/eKvfeKsfdP5lJNFd0cnVmjJ6e/dQ
PJYQXZ9l++RBjUgpS/E1HXN1m7U8Mzd6C2Vmw2hNyUajYMRXPhzWt6w8Z3trTkQaJH5xxiM1zurE
8hOq4ocn879JAm1REh+ZdKw/Y3IMhmzxFET/rt2d9las2V+rctU7GxZte5TgvLvZo2NCz8o3Gwmk
/XpAuZn6GIF7U82W2OcPPCbqDigmuebAb+u3D9ss3CxljqG9slUpLbDh8DlgNrCuOCemZ0GnL+Tl
NK03zQxT+BfVLAWYEBKa366TvSwrE7vPWz37AQh9ZjhNAEblvRuqo7ij1vDCK7RPQcKFghu/YfiM
s8BJ6RsC+afBrmwjIUGsgKQ8KM51sQiDMRSDSQOxNcXnMPoch8NSpmY4CTrxcgDC8YpNu3ApBxpp
0zyRL1igX3S3gMzI26B4TUDzX2U/R6DBdPoGbBMRJeUT592dOty+awXacJAA+y4meln1cJb2rfWb
ICE7KtA3alJwdLxDxcSTpthJjE6LZxlW+iucnsd4uMKkOeNToP7CaDnEsWwyhPwgDzN/554jQ9wt
zYSC8A0LATSOOJ+MGSjLukNbMs+vfyUXr686su6E6TZ+muXFtJIBBQ7eQWkpjNrh7r3uPybAeOx0
BS3EgcTH5xjm81ucNUNAk1i/T73UfrkWI6FpsSGV6jBzRuseCz2y7rwhFOJM+t1DmGRsPRozdTKp
FuxUx+fUpdxmuez0mENU9RP5PMPmDcY7Mse0ut/jPUPeR/aBczBuXdSh8Y8lPcayrr2IHpLLLp9l
QdA5BILCeCUEBh0ctoGr+O6BhaEfcte5br+eVqREr8w64qkmPxqkadrakhuBxxCr4nX4TKZqc1DZ
THZk+Hu8U77Zuj1L2mOuLdmCJ79An06vNRNKvK7C80BNTpSWyr1W6z5wH8Q9SipXCvB3mjxGRQeO
xpzJFu8dwO3IxtRjpPsNW0rwSQGA24bZCOD/DNsi+aKv/Dcy3Q5vl2u+q8Sw+8SE6amXBGsWhCfq
ZXESu+GyoRKd0JYn96HJRo3EjUd45Y+51pwPy7CF71aNlUOaurFouqtrAZypOr/ds+9HOoKDn/ga
0GwBlNRP1XsrISYtgPv2+ZYFy+AKhB2J7k3ui3wXdZwYAWkCwhI2gzPXlOGc3NDxBwnB34Uyk2mO
DX7I4BHhMTK93seyMKkbxJfdRhhi/F0m4DPInwyBsABgv1QvuIElBnDkajT9NaU2Qpyre0NaTQ5K
rFEjqAR6BBtc8x7vN525sO4xRYoZ2JJibSnKRR5HT1GJ7w93zN9deV69TB77GcW0HuzFjalIpdmI
0T4R3o/81PDtlyRcR7SDvgpnbQHLPM9LE32F0k/XC/LhS1QH1fhXZdFh7g1g1H3bRXhZDOG511Z+
5ii48wS0qxEzHF75iJLyOLqIUgiPAdaBbnZ/aayG0z6mZ6FJfFzZKtDgUvK8xOwgX+kFsL4+5DCw
AaZO9OY0qBJPKdzP6FTgYhLmiHAKroMtrTFXjS7GFqpdmv+avIfcKJFn9jycBEW3nJXJDMfYbnvX
3mjQck+0DSMS6j99uBoHuCPs9U8/UGkgXKhxTsYeoCrfJ0Jq0y6DD3WKI2X6DoG3Dd4OAtZZ4dC6
WrWHBz+vOInwzs3KW2FmofPIuSFM9JE+NfqFL46FS9GsAndRBXSIUs4QNpmpKmGwmPQorH8EfTIo
fyb+92rT1p6htzRvTVa31kxBoy0LXqJ+TMtN1+CzQ2u39kgR4xLySHsBm/iJwRDi1BxYZ+7g+CMm
y4nL4qEvtU+zvHGR1a463l2Zg2yyHa5cDd0i9SKz4XaCUhcvKoYMq4pN/v4+UhtSPSOjuDHlyrm8
sQ3F/mvP+ztYZSLSdqO7uhrLjDy1AEt0NQ2JFoB4Ibo8YV692KkyqJS8CyboKXK/tnqU+MKudAeM
evXEPJitGAPK7wTjpYOm5WM0ABWv7IQSgJkBJeEqXwx8YMIkN7NQBcbOIdd0lkVMfALx76R4X/oQ
UQP1o/R/UTi2YAboJhnwMiehl2X2ZC326UGJlin702Hl8wx120ro71INeMLNe+hQOCPliEYz90Ed
bT6epiRFuxRMwTXWu8++ur2mdlQGAEEkJ5WKyRgKEeyT1CrcP82eKnt/fDQEik1Up0U9Hd4g1nld
N6/e3EUbUFXr4f6/Le1OTrS5o339ZI1jjRtruHHgMamWLO+Gq9rNhZcfeyoIgYQbtTWFYJJlMJnu
GnLGvhhNyHXxgc/T4/X7jhGcS776syj+EqDNtEB5xA6lodGaFvDbbJEtHZubtUmlXLbtPStxrS1s
kW6KrwRtyPFiz9mrvbrrvnq2RJs0fyJeTzaycabDTwuWaMXCT0eiRBt3u56tbadx3b69Ap/KziIT
J6t/iAt6+2EGbsMZWNDKQDYCr96lBw9Grdzm55lM4IRkJRqC6LfG/5KfUa679PByQRXt7xeYQ9Jq
4Hk3pyfBIk0A4PtHUMAMSKdpSB6s9LlYjGyyMU+4i/tvjIniK4D3sjxlvv6XHUStqrKLOra+914C
d0LeVzEafp16WDZ08p9KPJp7ElJScL7ZMZ4k2wXGsAAtMa1VoyrRkTlTTqLC4QZwBjTQMzydGT9K
jtAjfdJrboTKoDUNrI3Ld75INA5AlUj6pOYrzkeVKptp9Hki0O6cgf0akB3EiTfKLAB471EU9CCk
HUTEC5J8fmb/25Ut4FPQqF2B3krdr3LGmBzYuKIE3ZrkyVQlmt1e9O7+FdPyitW/PlO8ZcvK16aO
LvgjlZd6eGUI+jm7l5GFwxSZhXZnWtfBaj7ltmXMujV1a5FwNcRZgRtL9/VOgCLw0VyAbqVbKIqN
isjv0QBA2nUUfSluFwxdQEyAZ9VviqmwY08zDirpOuyBHQcUBkvXKZMJRUnAk9CpIpVDAga0snbg
lq+13qqnM7dDutysmonKJ7KEDASnxYv5MWcBca6IreWU/UVnjUV2uxNl8RHn48j3CYms7+5x77Rz
eJCyrb4KtPyZySktbyewTFKRNTVK3B2bp7GbmF3ooIhsZo9v+BX44QYjsicwwFMO5DRu6BLkNSbq
FX+f0PGZXIYp//qmpcc4d5vIG+eiNO41+9c08fzz8VACfw4IPauF26q2KTg9l8RZ3zeNuUxmrmEy
DMYusLLNcJZbZMe0Ma2sBT8+yxGe3z7kUqvDzZZdoOTrJ/NJ9o/Rj1W5xJhVADHv8/HiHrFzsQma
nk8XNKL+u0kEjN8+EN2DVaO3abqLRBmi5KTqXUJVusv8TnZheD1BFM2M9rJ2k1Sq+/THY5s8B1Uy
qUcJE8g0pheH1R5YzASNOamyGWQm10wFxt2uzXbeza/NcTymU2XAzKCvkWEWBvOPFg4UpnKqyaja
EiAcX8feD1SbM7Tuw933JYgnGiaMLxJbRSLuMd7qJTnQgj6IdIhKfBBjPyE93eXUfqCp306QZrhx
aUExY4Q02btcM4ehM4LbHsW3jNlXkGmgr4+86DxHi51rPjUWEoMuFCUNUR10+IibA45n/IoToBYC
vaSbdJ4AUnEHb+8lqJaSAzqrMvZAAi31Vc+Ie5Mb90dNvvi45s2AVQt6f8SzfOYrWbgXzEPV6DwG
rOpf5qDKU8hYC8mo8xrVgsUVTZITEYQkSzKjq/gOa3CYdz0xMnDaptKABnIBM8K/JY/PPl5xPsx7
7SepSQHjShOBmRKihDvNea72B6SCvDRdiMoDrJQggHqNHSwCEIIgZ3y795OWURyPLnhqTTSYEcYt
HVQ1d7P0IAMaIwsIBqMsBHY2LO2ZhE0E2mpxebgTH4mqQrj/W858aLJMbLejUuXt50m3GlNrMAoc
2DFmUHFnJd3PmmwVuSFzPmCzh2TjGXSI+DsU1RjYguTsr9oZKcAUIi7F0F7v9ezQbypnL/Geq97f
rjQgc6jFoTZ/JoraThsgCvCJUoJYPNlslkY7n9vJ7BeLI678bER38nv1o58VRhefWAMNkqkNKbtT
8r1spcvAqHMkE6YAzAvgAJ/p+nXVGx5t/A3glgd8mWwMY2p/p4b89qpdw0cofFjihCUYFbOsMcI1
SF4+Mx6N9FeR4Gn2smoJWl2TUDwQcubkxqanPc94ugHovXFub/soNbg5ZJQoIlfAtxFEhReh7Lt2
H6p8X+hdcJtdN+IgUv0dXHgBjpLU5LCi29d11YmNflXppjyNih0ugEUqTOGEpI82fFPReM3Wwaxf
GraMhT2CTf6FZTybEaVxSTQZNtHb7FY90bHrn4elSTfM8AmDDZKZpFWCVzE4fi5QISVg6nXEsPks
GOdBvTmzoaVASBps7biIZHoH9/LMafa2VxYp+IVyvaXxqEBzSyfMREgrFrFAT1L+3f4X6F36Bpkr
kfXwFsQSK6+fHO1pWSE1tmgKJZE8ag0lmv3+GET0Gwvhk7wqJ9ccllFeAhh8fnpACqRpK8a85v/H
fIAWGcI0b/6zrzcENGgCvKB/x8In53rkoHmnWdlm3ISibqz5ivclPcQp201Xw5GXRJyR8M8R0gAD
RVVteE60P9anlojtpDQEc3uUPs7Kq82kmUNalH99h8ZoLGwAWFA1qXXibDQ1bFuBh6byeHRvDOux
8Q9EdRFr9nOhLEFiaNQb8S6Re7CrHSjsXi5aF32qB3WgxJHD7mtx2J9hns17OwE0DbRJWgBpfRzV
VDwNL8OTATGZSJkgefC3Nukca3yBwwgfxK5MWXpkZrAf0LOl+RTUr8ntEeJfdrn0rf9QzljW5Pvc
9jZCWrf+CsgjsNRhPakss1PR5HGwVYbsqPRx/1T7ii14ACVamo8KiD8Mqfc7pIKHSpNTFzzdSi9v
vA5R/LvN92f9L6nHFp0wkZTz+5NDwNcPxf3XtrHRaU/EdUvSe2qyuphhn2t7dbkaHx4Wc61z402B
8yyjm/cVsSAf8oNgr4N6InzWdkNBHUF6RUQA++3uUVQWEMg7UjHc1oGe1tYWBEh3kNS3bRGPAyAu
nkORHUVVV3htLUq+RqmqTZgEhqE9wBfTGEgIwX//Z3AGA8aGft6mPkRW2xpIBYAAcl8FkVycE52G
Hi7RqiupiNxtMr4nMYGCCO1U+vHlVGKzKPywEgH6y8GJ6GoEvHnvN5l2q1de+wK6bkm4HcUfppY/
4mV/C8lf2oGjSg0anwEFF1MTbGeDNFcRoCNKbkGmGnAd2s7fuQAjs335JHd39+SFNTFXZ1YCQvqn
bozeFvH2NcbdPVQdbK4tQqUDQJ771JhfhBPDeen7hr+/SgMo5ZRu+CTuGx51WWESLGyVItu4sxJ1
uSzV4K4PiufCCHSki+vn5l+ePUvHvibiJ08ocX1xliM2ROCrNgLMtEO4DovbYoow5BmCMvMK454C
rpjPTmmYtRJvCL1gmYaNyHl8/3RiEY5Gosd22eAWcYb4mpe+jT9+NGS1e2yyT/4vNwjYOpTcJqiY
9xqx3nCa7Ndwj5dzspn7Rqom1vo9H1MyX4zViUUsqiXDr6qLI6ESnYybAuGP5+xpcmVFUZf5bxK4
Xp1lPk37+umm6itVewAMOgkoUg6wfmUxhZogsglRRjh/5JwROSouobQ7WxzNlhyny4c/ed8/nX6p
eZfXYJPFllCkkD7tLvQzgtR1uan4GMZGHcf2EtGD7B6bPP1mUV53NABGOoesZALZI22S28fss1tT
IfgD/SwQKn3SvjZYPihL/vQg5ZRK5fkNOHuFu5YFVx8ijiRwbVTGmNehB7s1NsjLDEZFR+ZIbbhe
0WZEmQRnVMF5TxqCC1UMwayoIaJtDjCYMkCAscKp6DiqdxDHXt4+qLVRgAmKP3ZeHRXYnKb+6Ijh
vxi7DxsBhyQUGw0wfp8hlA27JTOS9S2CwpOxi4sG76jmyWoPF7bfoqdnroeN2ZjdoynXwEa46ttr
PKjCscNvgdI/nBmU+d/SFJjEqLAGNf9ZTNXQ5lf3ULZL/YBe0iVSKjOq+58hnmg6k4+DYny5lpvg
CsO/JnmY//B7q+o7qcc0LbDfnwM0r7txzn25G5/GNYonmPoJBRp2vqrVAtpqlpa76dBq22Xxx4FA
rXXLBz54TiZvORZjsZ06cuwoTCNmG+psRuJoVOYuQxRUQERuWPGHHVbQ9MZAWdllYJ6TpN2yYQVy
lhbJe7uA9s4TYE7AX9veKtu642dXsc0jDz5HJMHShJ4mecAOvX/yWoNCIMZRl81RnL7yx8n0uNu8
x4CKu7T19uTzC5q3i+BtjBR9Z0NkHLv7FP9nK3eLg75uZ9fwn0Cb63nVIvwBx59deGV67ial5043
LPHxusFL9CiANfy1C3b+gk8vwQYVnqpNCI1lEHCCT+pPZlnrOmBovvXogHYSlZ/xVqPkOmwDESOk
pdQ8OJ/baMh3R3WRqiOas7S3jVUyw7Ygdvtz1HG+dvJZ9BW8p58h0gQnKbwNxH+5IslX5Bpj8OWC
7uelfppevLMRYaXwpvV4Il5R21q2hEyOpZNOjHl6B9Sw32zNNQwz3dfZ3DD6lWlCXKSu1/ssAPdp
P1VFYUXkXiWyjaevXeOYRehIi/6QjrerGf4ujymr82idoOmiPMK3NNid5bAlZ3yxisEjX6x1Jm6P
evN2fRUH1Rz6IdWISJ806dN2tEbM+C+JN4JEIrMWBfTlgysG4JAuzgEIEgLBFvu3holVuJ4/KfnT
joz+g/dzZ2ciYWUEvXSZ17DSEou4lK9wG9lPkPEDxwU4IrfYq4LPN0xSp01OpkCtZJSkRd1I910n
NSzykQ1pXdfdpVsB/gDwpvBXX+5m5wHOYOovjJeumIMr+G+l3nxdNkYqqCaIngQO/jc4Eti7NdZM
ViLHYvGMpLEO782oOUeI60xUOiraP4b/KIraqXMaVP26eK5VmabWilLKBlX2k/95esm4q+dBk62Y
J6mZ2SKrilGp0VBdG6Vg4Bgyo1ICcPdZtr7M/KWepPr63e4/naNSaciwO3P/1qcHGzEYdtI1LSH2
UXtcPxoyvKqVxu1p8T3QLk6eojTP0UEtJ8NYV1YKmJfwc4SeQYgFOKxg7RhRLevyaHXaU0bTivGa
1aun0q+gnGbymtA/0hqBDL19ntxdWuSIqaaZlprzikorr5Q1GyLZa3C2xhjAAddXGg9nd/NNaU9C
4uEoOWGaKw+YpmNY3Y91znfHXlN+ytkaLOuisGulScymQs+ztgahEQ/Ki8iu2sZcQhrGud1V3qjT
8mytc//Qkc2Elqhx8ryP821qTKjbmcquMTF6rQXlbBWbsVPkZ7QIswHglxKfDeefgDOBYb+ebtP1
ytswyb9mG5GQ65iJXz0mOSLf2PZlLkVtWlYQaq4JxSeQmz9F8KUVhVDDfvNGF8At8QxXbVJ147e3
Xl1g/3v32YFD9YOYG3g0YVl07Mkx7i6uIkpiE3VVrYN8twJ7PpHBd0B7uOlJ50XEXIsykEJh53VT
xLor2YAfXtWVmr06+1lqAkzNp+3vyNO2F5qS1/RfFCTuLBKdagZsfEGc02CLLh6RsNrM40DbPpz9
yH1Mk5KSd0yY0iqeqTFxlFq1mifyWdhfMN67RnVEWj0sKtPfsGQsCgnkZURtoi7zWpQ1oT3idHlW
ndZat1V+vCctBa80Y6eIcmYguxAFC0ULS0WlrQvaIiLZ6vOZgFx8Js7Lkucs8QATeLksnl32ofl5
cRt+/ytPqXhmxj2KLUZQuzwsuXMEcbzxZxcRtAdyFjhQAvErYdOlveYB/hkiA6bBu+oAm3OSMa6L
wr3gyzLICRmvyShcDAAOsTBPXVCafowUxCI2S6gCCTWHQBiWKs/wwh7I6wYMt5jZDyyVx6bmlTbm
Ai+UFzSDRENAc2GTUT/VRwCN6IU+1W6ORgbtaFTZyi4VKcgnskFvd4xIy9ggLzQvRYuoDA2xXDRE
PwGtpJBT4VoFktyiyG+lvz4+qyJBnro5xJFZUOx5jzfUOl+l2iisdjZeMMFFrCi6IG67v+OzSejl
1Wt8LHpvL3Cl/A5eCB2XNtx/IbjrGTKuAumoqUBHHRwyntDp0HRr7PQXMQg5qIUzECCdXDKB7zLw
8MDBl0esyfGqk5sfAxm0UaBiT2Yrr3iB2kB3qprnCU4c5FSl1msNI8GEplxVMSebB7LOvaU0k9dO
xU3R8P+8VRFao3FFNyLAqbpzRFL+UQhCfpe+2Ro7OnnHNaK4/XavCS6aQA6ozIlnUEgmDpqLFQpm
ZayohxmZAluAhB4QqyS/d8JOXGyq66z35c9Yau8SBZKbFiXDuwh1sXT2a8ghBNlvGU7IdjEFGXAZ
YTrUQGlmnnHZDuIxL4UcEhLlkQ4QPil/CunY2pCjcQqS/7nNJfXBICPn8r9lGIi/akAoipq4bsfp
geXFesRCezAyuMm9+96akhJ8z8+/ERf+rKz4ReM8fLnUrA/5exO7eSe7cErfRFe13pf62WCYx4Ni
PLggSQ2OHmbBJ4lY/olkRGbkAaEaQSZlmMZVw3xwRkwMXbdfAF9mjbqmHF89TOED/Fm4Y7CXS0C9
4iiOVMdXz+eLs8T2o1rMbvEZRg2fuIBrF0QI5R2cRfo9iW1kB/bvvujm79IKbBSDs134cJeAO945
nw+mPAddhob+kJaOOxtMZalvv46YF0TrAGOAu0EQdxPZjQMWxMIAcFT9D572oT+F/NqiSW/2klac
9/eVfZ/Wl9xNW2Frg5uDyOayT8PHMES0JtN93AT7evqbxzIlMTDSjx1UQ9CHMrNy3P7GeegpVF2j
apz7iSIGIsYZ5SmWgJ8XjqagjmJNzRWiDkYxdRNyVbrdZ1jjDNoutEL8VzS4Hi0E2N4+tP6tPyDz
FF+/RUVYB9EChbYPqQZR8gtG+xYohhGrw7rXPjvlweC1xq3uwUISpyIndsQQRAQYotiLLN/Yq4IR
HY3E5YeVAhmih6i+eDY9h4WNR02L7b6YynSmcPzZIa4IpJipEZcHABUcdmOseXfxExgHlqI9PXsk
uNOvDlvG5zCXmJouElmuexs6lyCuMpxG89HG6PZ2+c/6Bl8zCe1IpTw/JU+3FqrlDEgZKdnLmkJT
0jk/c8MkomHcz07nXCyjMd/MyZ0nwuB72upQOIppfquAmDeaAP8VAuaGU354tu8QfWV+BH99OseH
K0+F/+fO0ggvDG2vzPmj7AL9DB/PqepppmffyJYOJbh1pc6dTVdhM+ZZXNjgmz8o+Lfvf1H+Q8TO
rgIImx5kBD9HiFWjHKwtKeyFNqcjZ7qa0b/ezBC6/7/gGU6VMnxtlbxAhMcxFZByGpsldM7c71ZW
OpyJLbULpq3tOjh411MEKAC2lVLZqtQFN5gJZe0pB6ymeuRg2eATu3TOz4EGI/LHF6hkP/bf+jab
m9j67DfHvRF61b+owiJnT+gGnhaV6WYO+Oa9XB9HLIzs7anSp3rbP0kxsvZ4Bpra+benENuSYvgR
8t339zE4KgxHTVmFbdK+iCEN3uPPI4HSgAqpr4SLlpcNE0x8rNjyGrGf8bBnXKhk0MaMYFbAGGVD
Gw4dbmTfvn1x9cW0wPbqSNYNh1lXTM5ILRio30CZEDKWCRLS0L7Ef1SO0Lh/z3dFlBDPpn1ko/yG
0pONT5TAMBs6qDMBdngdF5mhrnLKMVJKT3Ud5YxRYC0Y9LvTzPVeblYZHmbpF3lRrT3DCDIMUHak
ntTN2y4jNW494rWy4GcRddXnHDWLpWsLPTPtNH0TUk/qQ3HqzCH3fe80mkzgji7/Lf2fmFa2RPkK
ckm8fNhO7AA4O+7g1uSiy2o0ScR6FhSpAKMeU/BNs8n7xfGLLRq4aVMrFfDBgqdneYFbheyriwwD
BeLPylX/ATYznMC/2VYleP5aC7KOsasPuNehcsIbyatkjMu7uEnbROTfq2LlAavYppWRS5yvfUlU
LSjNQJ2b4YrQ1uMfnsQaUXq9H9EzThuRmuGUDKvrP8XxA7HXru8+zfWIpBCTEG/cnWVXMsBn2Hcn
VZrBr6svWrWUhb4TElQM7Elfi5LL0S0z4PwV4VvlECCs5/djtrtWymoXVFDA7LxkVhwXS7FzY9do
vh/g9IN8+1HiCxJeMPPcvAvgiXdItTDLu8GEGlUEsOuykNVNZ368grcXJoTLQ38B1kBFD/Nlvfzs
amDJ/kGVB03ExxoH8Eil0JDbee4tBGASQtfSTlUucixkI5gxAOY6L7+M1bUmi6P9MxYNUWqN/rIJ
aaYx3zMb6rOTLk8hyGFsxOLauQYwet5xGbz2Ql7BQyaoNb0bj0+OBh0uBkjEqmsNaYQasoRINeIj
oEUMsNVpAJBeNy7qcEU/ZSGDou2x0EfreG2noBP3eORA+ypUVdxyQ4rPq2Gdgg94ZwhFi74tVS6T
/tPmLEHHh5tZm4KN3NgesFwG4MhPOcnkayQlB8tsi9EyYu6HDZojtXwPL1cir5n67LL6yEGbmCvM
yTXob8a1LkczThbayFgmZpMIT40+evMf5EpCCibBkrj0bmYR8Gv4Kpkp/5GWYGkgDH4pHm8K6MI7
UtGrU7T8g/vszORwC7U6Woo1Y4pcTsJDxiCbAN0nggXHnJlIhpF3SBGls1Z6tKeN8bM4jvoOdqLI
68cXT+h5+SRLKM8TD/XTUmHR2paSFs3g20Mjig9p3CKXTcvLJSkBdHkgUKQ0UUXPQpd50Hk6uDvu
M6SK1JTV1h2xLdGec+SaK6ArgD/jbwOtGjaVv1+nNMuwq0o03d6J09bfQaEsHXYk2XPzMjJKQH3G
el/xhSX6Yf7kF+6E8e5FW8qKk5gZm//PxNWtZ/LCABjUkqBiL4eue1zNhjXlJmyham41irK1uHXY
Yzur3rTThSElipmmbr+22uA6m5VArVIf8DLvnAcg7M3rZOMMUhfL1tYb1IawK6+3XvwA5mbM7yUO
l/2hyg+tpi/DDhV6jNrEEgU/CCZYyDWCdKdnksuwM3jRlXYF0W2i2dT6yOqjYhZnfSWtsn745XSQ
twYuqL7OY5mvGTQo/T2r6FS+48AkD7Z2wATz8haW5mmaq1mJgyZUz5njazGt2729vhJBmuMooI2s
vVzeVSk6mekRQmAXX41ndfc9ae86QgbE+fJM80uOX9nSGBGX5PI/j5ShXL0BD+6aw+AurbBCNXgt
POmpNObMgJi273CcJsY6lpTN5op+AGgajC8O670tmUbhB0cM3BprN+ptglh+A3xCNB8AyQjo2mYF
983/zWkoryx9rY157cSTGAkRMX7vs9duKCjSc1KsW/0NA+R3VrbWhKsMLsbGu4VK7H/dyndC6tR8
YacYkc51ob67Zf2KnvRhikO7BSWet/2vlo5PU8Cx2RWB+FZqGq+u3ljAplEUYIN/OophIoMDs7F7
L1qH4utcD8E4IpOGU6j1QG2PR2PTmkRTYPDmKe2Qh/PeBXU85Dv9wetuk/hwathKnjBsI0Y2AyAN
viMFugOs6D5uYuR+mGzbtRPqSeGf2zEmy7U4H26ZqfIMcPeS443P2pYXuLYHL1vaHlzwM7QRkZHZ
0Nh9V3fjxqJOredbfQGs5V5XgxGgib2EgZFQYTJcTdXgHYVswxTcSwRs5Hll/XdvgNFFIjEKEsm3
Cn4y8aYdPYrL2y4MtE4pEGop6kFliOkbjMttvgWhPqfsUNxOjbG0oZGD0NwDWNzFsrKQos8c2QGg
X78dT/mw9F4O/wrDgRgq0L2hRuC7K0D/kc2J13Xn5rBJSK3dkiL7IpoNvU3X7LbvKlc4pmh7KmXj
B9BIUikzTXuZepBDHcc1sf9AgPgChxaPFa7J3zpXYu1kkmV75pzY4V3DYP2q8NifkxnAZnJ5nMkK
OreSSRMMc+t/KVGX1gXZ6kO7C3dCdAQK2Js9gC5U68jI1bd9f5jbODMTPKuHxwaI/ImTsImL8EUv
0hlxDiD8fjvJnBWnjTF9D2h/mxQrmqAobdhH4RA+iNDxSdDl9BkD6+6djy5PEieb8wWRk6vgCYig
xPUlgBC9ENxI5Ap2FyvupXmJTgUgX2Z7RVw9KaQojhbLlwnTQxhySy9xes7fQqH+s9gyQkYB6Rif
KH8OVcY1VUSLRG9Q/0PLFojFUqrNhzNDO6D2K7KYsYp6HTUroU43wQi8UuNoFH5SWh1KAhlsJjWo
AegGO21MnZvYdt58teztJXN9MlKICNgkRfuSYRNEMjk6lRl7nWnV6Cfu9Ywev6sZIZ16yg/kez8z
lXroZLhZuxfx2XfOhUQtQDLE06ayZ8JoLnJbcKaYXki9NDXEkemJNgJe2hc8qvLHXnAmwJrNXJ9/
zxvOLurR8bHrfhNoHaAcQaYO/Sd3sddnhCghVzbBX+PqwA5BubeolNS7OFhxUCHpTH3GrhKwgPSB
btf969BOb6yRDbAcu84yCEBL+UHr4lmxomb/HhDRdjfLLYXR4nM29IVl+xttREUbgAl8qigmOPL4
Q5URoFPqnrqIaHwPKB67oO0mC//my5y+H22ACxlcTAM8hPLflkvW0hRvvCWmCnuqTC2sGyfPlUII
amZ87gOo0gzbyq57rSdReVYgwbOtwSfX/qk/44N2S4iplqS8wkdcAeBZUXNW4eOafkncHZFXfrm3
S3QL/ehVQ+PRAohjc9HPOlm4rkHbSJihYBluMxEUsPGKrV9fzGIQ1x/a7C19dhw898dVhLf9wWWp
RBZqYVKqgpRB/nVzF7RBJ4eekhIVEAIxJHkgk/Qz6YcNuMQWWn0u4d7zJVE29tR7TYG35e71QXsV
tk47XwJvuuF2dCNTFj2eKGImI21uYxydfVhUZ5SjKfeSg7mRkcxPVd7tTG0n9IsBkD4iXvP7Ij6U
QSXHIghJL0T+C+6NC6K4gZF9pm1wXk/pJS9AP0mSZxs9MKCjSGeiONSqhaInbdJxYDjFBwy0HnzG
mE88xTXTyBTtCMa5P5CesYVmTSFuNmxQCyWYGnmbBNhzIHQdQSB8lb69e9XNtFAGoYnFw2LPuKdt
nPDUdBR7vjRF/iRqNUsL/kvzeLrU06sldoH7mizHF4g9CJlC2pczV8+C2gfGukYUXIDFepsKmftM
T+GPv3XbEcPZIJK40R3hGpT5iLCE5W+5SGAnL2Q7hQqq1RWZsT1q6xG0YcYFwNdHK9FQ85XX11yc
uZn+oePOpOqG124VibqeudmbkQ6UlZlEjyFckzRQ/N/Xxfz5Fre3xXvoXiR1sE6Kb18Qy8fowd8t
GVwvIG+bpFuIWq+Rz6ocvGkhGkO9ClbGoLl7vQcLsCIsDFkITzKhlMGFIm+cP3uVks34YJV6mxbI
IOGNNDkZCfJkVv1yQ5Pe/yxIu0EJ0ynsVSrFERX4+ahEdkp62czpTiZRcTdR+gKfjwtwNa7h+VLm
KSvFJy179sdylL6zK/vkefgxRQTPEA0G8BaXLiEOC6sIdTHzvMN5AQRPg6s10C4TRSx6NoUVL/Rg
hoUf4udi17iZ0MR5Aiok/OMbyVJl2ehraNeSNeDUBtI8l9u+7SBAy94TQpmaSRmTzupbKqpf0O2k
TJvtiMbE2gAIuh51gaDnJidOT2dGjdu4UVHY2PaTB229WZkC9dSG+kXhlJwNv7EUXJMcChJGrIMC
1GVtyY1oW9gZlbNf7VcDfciLKCuYfUElkZ5VdVPv8NSrspSO1xxLAYy5knUKEFaIQk5+UaznZTXO
j/HnxUfApKEyq+0fNI+HkGNPcdPuFWQrAVo67FUnSJim5mqIQRg0z+usSJYpeuKX66v/vz/pChF+
4y2wa8y7p28vbp9OzV1nUXViDrFh467z7aWhxP/cKe6Wfxde4P/uXFcs0ljWB863M1cTEc9D8uq6
iR3W+1ARRo1f/DQWBj2U8YufJMi00mEH9rIEv/Nw/3GfFiH7ul6garQzZbdFt00tPET2C8OF/gnZ
NddNLhj4/X5BL1qGLPycU2kBlPSGHlS2KjvEIAs0xD5LJiPT/gFIxXpBDmXF09H7MzztnKFsEBHl
Rc1jsryyLLUaAlqLlm1noaJO92s/z7zHeWCG+gt1IvoqQVoAqGvCwMRwLWp55jwsJ4uQ0lZiP2S0
kFMQKS8WmZC6mvtdG2nO+RupEdZHDGx5nWpcQM2CBZ1buAIpkc9svrwsXQXtm9BYwclJ5QHUKLmE
pV7T0BINVzuOudpiq3jUDs9fBDJFPpeVCnLo2fwLTQvhtEow/fICY1KrZ09qbREGZryYXlxeV982
qbrSVcOafVBGHqYJ897P0nwRLGWKz16EU15kVe+yg8P10UFpQSaqibZSonJDdIYeKZ62f8y84LUb
Kws3NeLWCVgqoO9eUhOruX+zpnvR9IHaE4e19+rw/MO4ST7hxb6vjIetXS8TRCuN76TM3M/WlIlx
DNXyMEfO93gDH9xnjq359+e/R5FVBSLWNFfKwbAKNfHqnl0qmrxTf7naB9QTafvtHRd9PjORQhNv
RzFSGi+eZNxrCvqaEflZsKuvMa1nCQ+aQquXQKbHHhrVbm6mOlWK3Up0mVd2izUpmGhgEG/Yihr2
SFMp0HZIcta5wa8yy1MWX316Vl9FhGniXO9/TH5xZatJ6e8DVceIVK5Dk1rvbP3cJjtAF9JDlM0c
fi9NwmXdw7HLNzuAshN0naozs8GktCkyxDWsZmDdbMyDQZPcFw+xYkEWGNJy5L3ncs00zlWIYeG6
T3RNf5Zu8c3P/bN3GVdcEcUAc07o2jnhv4QESlparqqn1fRG9TeWBC657/5bL6CuEJ5b4PAjB49m
Ygen0zKQXbd/t1ISyUzmYJXTn3PVI/FnlmUPd7yY+y3Bx+H35cwQhS2AowPeOw45i/zIkA89xlN6
Qm/oaJygazHvOViIkimI+1UbxLx+eMvtjlqUi079TrLQJS7U3sCRGUdBvsM5FV+c6yq3fpeA8Mc2
8tndtD6h4J9J1i6fkAtqxmI89YRUuNNZKtxeYJDPEo8laZIYX/F+8Q8glwSU4Mup1sRfZm4oCrFA
hKlAmm10nG+jvyQviV2Q3YOLQDwx0WRbCUYe1bJYar4yyu872s2cBguWUF9BqDrBGuo2Z29OT/B/
MrueB6w/abINCSiqwZpgibQ1hDVrF9mP8DZyyaiNbkl/eYkfQgy+skUDoZplevLWJmJv1j3EJz+W
jeFNyT3PgNqLB+KtApmNvaVVac4MZd89tC17JyngoyDMV8km1j8IwSUoZ62mjSaPPfucrPiv51B7
yGWvvKP2FcN+MGQHRu2rnXtgwG8YJ7TFVb84k60+kJVYM0MGAteHBazRK2HfG97xdn/+Bdrl3cL4
nsnY/oWxWxoxDaVivenwtGqHLOLYz4kpFCzITDqSUGelwoxPLNoqx7NwiOoC4lXRTNWKJ6I9pTaV
PT7HcCgLc04fyQawtj2aDpRfefLK0Mvetii+oOGS+cdk9S9blnuY6zKgx3Xyv17qFDbZsgGT03TE
ZVeU3zQe8Q2Ar9SfBXP5aVrnw3ySyNDQSyyXuJh1yPDGroU4Hb0pE9VdlgASPemMw1YtjMd4AA1+
qF7v6ur6MEfo8uARc7rRpXUAzwBNSrgrIIKNDJl370tvxmMVhZQ/deldpcQhxyBUtpuQx+Epe9TQ
mqN254vszZyQiq8anB3L3gMWT4cTMtNsQTvT4+WdpR1LkhQaQumsu1VqOL2I5Jw78alrIA0FtxcI
dRKMFPUAy/4Ku7kFFTba1XWF/hGaJAWttBLKrGcUboCqePbuGKViIUBNw3QxwbKv8lBNOZ/RfxJK
/piKr4RmPWKluY2VOiyW54sBbVNgGmhnL8sTK2buWV3W1aOhw6J9xmGYcSMh1nrT2rzHntV5mISC
csBrcfGNj7eSA61E3uT9qNFbIFyKEtwugIBjDiLO2aja2ZC9V04rwB+3/5Q7jefsrcHMZkBoTuUE
AwQc190JTzYLGZzfVN65TpiETKn6T3u5TaA1dyAjbXzQKA1K974/Q3TV8iwuLCpqB8mf2c3/nTjh
1+Y49/NT/crQ9updFbcr0OXH8Qeqp63BNuloVCitLYWzCVGMkEeXf8Xu0VHfjjhEf4b1XaEI7uwa
lAXzkukWXWSIwZzEU+hauYh1gany5luSKkR0VRBJkYSO+Z9jTW7RrwLpmxunumal+orH49mytqQt
HBkNWd/SqPQ2QpdI3RGyXo4spOsxT4VrsBDCfSO0CxQmq+hz/1Mu8GIG68dfqF2dYe4kf31Lt4hl
hXJTgFmUna6Qm6nUAkLDQ5NwV6+5pfcFvSZqYY4gkj5AXaRqrMYNHvH+E9LnUBdIA+6WcH0RDAOC
nxR3cq9YC0VVAcnwsrT2/pGkljmt6I64LkFiArkXs5JRH1juyksqxRpbR6iOjkzlTXcYnMdPJB1x
PyNROFW5jLTV/wSey7MVlM0PpwbVqvoT6rMb5HZmXNATpmWXWD2jdNwbL+DDLEiVODu+ODpYgr6O
+TF55GYmYWwsDC7v37INOFxwIl2KnV/GSLjNl4kpIzVWObARsR/0r8OUff419iRmPNLG3vOLM2gU
TFdf3lu2VcIE+Fp5ilm3oxSaONTovEe97lvPT8sSbTsKO8MS0lhwOSpNMGnz/FyG3F/g28N1OXPH
rO5ZsJGMuQqvUeTmv8NgCDA3xAbF4zFI5JQ5zOYqRpu9EKfkAmIOsJ+1duOI8YH+Is/kbNLcnTn3
LUEw2XFi3hjm+bBdA2G981nkcMQDEs4zFF6DxmjRHKSU/rQwJruxJes2N25goczOCvCXZuMoYBja
/FrvKaF26cUAkd1U4W4xbIM0IAZ6tccBMJwMjb5wBR56GSJ+FJlEIsuyDarbrkCGU8mrnuIzxsrt
L+N+kLTtd4t7I88gMowZXovaBBntvxxvibd9OlF8rxVsqKxUpaKkOZ/EIZJoU23GaGOdWQilKQHA
bEF4HI21LjP86wn/hEh7nFatr6MwkGw4vJZWHNvGnNH5/e1rNuYjJk0dn6YGecLdxdgtn7iH8ygY
JmN5mc2cVYk2yKScZln6E8NnsOxtvoqbrDAh4lmk4oJCS2dQdHkrbXZxGtxcIxnw/ovT0F/HyHHA
4K81fE2hAm0G0lKIVZ/r3JdOxBZYjmcydl1OddhTUJRCrELiVeAZMr5YgRtbwXbtef4ckzUlwudN
UMjSXrkLKDab2KbUpXaGIv3rE+j+Uxwxkmg4huOY4zeOpbEXd2fQ4h7QIvrMfi2Dw/aD39N+u9JV
LfQYf5nJboZc7FG/lZTDl8yLrZ9S6rYoM8kAu4fV8p4jml7I5Rg1x7tCGLgiD2my6Iq1gm5e4Ovv
yossXuNv/BUORQo+msgHKYjgRpljjVd6P0VWwikpENvQ0QjYNt6fMHp7N1hUIBCGNEWypn9W6hIK
N51UTcibFha5yhTd/iIqnKdwePNK5EiLMi3WIXfYCAtLUYdB+LEIthv91lBJ2YeuhQn+9BfFAHDy
5gG9TTw4CJtG7K2WU9iQvJBGWQ9vI+I4MLVzEfIp+55xddhVRsdtTWlErMCPjXW2x/9cwfD+OO9E
le5u7zlyrBxGtYD3LzuO07qY6MJiOFYVYXASK4qtSlLYXxJ2KAeJZUfDnHZk9Xcsxt25sVy9ETFC
GCT5onc/hsabLo8a8tCbwJ6krN2VZRufwENHi105LlkpNsPlgXTsKnKT4Zu9+YYDew6FCc1bQOWu
FDb/BwHxyZfXObXjoNYbujGYGlCLcU4mVBOq00LZy4a274x2L4JYwVtQaF9Fs0nVI2rybucMNl+1
2/49e5XkWti6lHzkfXUhlGje8+vgTrcGeJvb0C5SuTxBKj2W5o9V30RMy9htDUqSuq60XPoJ3yW1
4hh9UWAqSchI4ectlm5aDcFFes5/WK5YuzCNC9eyKZF48Jy7skgJwwOI2O9kruC2WbCS42Ie43IL
2e/LxtHNdi+zqC4w8AhF70HFKWJOwDuYgmBRbK5xNqE2bSYd8BltnnmeLAfyOacwX72QDwhxTnyE
t/tWehU1ojfJjtYGi6wJm9MqzRKGshZR9VcQuKhBn2tw2yj/VfuO5IJhEwNb1/2NTEhUURhpDx04
iwiiAJI+jALVYUFKmlP3FonUQ/yWo1YjJ4MATIMYNLMWtQ7LojBwn2hP4hd7SkqAfERNs+rhSrkm
LVI42vkzQBXjy0XQOKOiuAb7GIYPsH80cpbZLFk0iOGKrueE5T7o3UGi2XtiXGDX7t/b0PJIQSfe
fAJ/jcSRHfulr5zJMxST9Yo5dLGXSVNDOfN3sh/G92Ki23QlFWDRNCDbdCHGidxn9j+z0EP3nuHT
4ZSnH0McMEF54b3lqBq+K2ea9q01OyQGlDcp8I7MSZPwFLZoAm3uFvXRfRsrGiNBcR1feoBXSgpL
UFvd4XuXbObe98ak1pAqKdG9HUyBawd0AkJAbedeId1Fj2w2AmdnkqvMbdiOy4/6ZLZMjNgd6oCJ
dRmytsCFLowQsX4hV1nkOvEyC8Rr23C7YMktvOpb7HJphF4dJ3Kak5q7NCBGk/jXQQH123vuUZPG
pDN8bqu1Oc/I3KzmkZDOuO/AuzlRSmchX+ZQKC0gu0GDgH75bi1WoVQk0GK34IdPq7GggUuh6hW4
i9ykd39VSL/FtqiGKZ0iuLa2ljT5av/uN09YBf+kk9n0gU8/ypUR5cm5i1FS5Yex+xV4d8iSZvuf
MWo2j9EOluVNwkorwXAULGl2BIGTdRybscuE87DwXnVdngVSMErGetPZwgoEUMgcGKtZ9RdBJoSn
bfEPZQYqhZU5w+OYL+aT6xwwVKLJl8hdXYTRann5QBdqi229jSmtG+jbEpSJ4oQU3ATIcBx9e8md
3S3glV82a1VJmfzvtxU+VWpA3wQlZGwyI8W+2CZfhl5w3iokGhSzHMdqewx/M0nsJtBdBQVjy4gl
v7sUX5wE1Q4KjCtdHrTB53ZFkPZI8rsNEXnePVOJq/2zgeBSobTKOVjgTcGwCr2I8Ra0xyy6KzDM
R2MGmvkSNA54iEh/off2oNUFZnnPA0XMRiFoCOSVdi7lINTHElDnkTOpjTMBmPtCJ7N645I4hyDY
t8ltkDqaTCYqlqR2zdGdNdKDazwUoSQoXAIxJwAB9f7mRu1VC9vuJRpurkiXyHXvn3bO5Yvl9a4o
4Ob5Gn0kdRhVrchqL7QCdiH+S8tGXBtFzy6oZYJIGpiSIXqRqG7SXj9gFgipwEcpKda0JY22nL53
jueQz7t7CNMzqE7LIBpk2wJ1TkHelQiVEB0uzYjHBlcmc8+TzKS18LUyqSbj+4JH7H29bexR10Kl
Gz3/2ZzIEGO84qwBGvtbDq0bb1Nk7QlhfuQxKcJh2kNPvAiq2/uBC9NMHgJcCMoxjOUgZlPCd9Zq
47OS+/yKT6+rZoYYQnAjOYMCua0+0aW2uVXIAby4OEYYpRWbj8qkzGP8Sc8SyqDMtVYHJhfQtegJ
iKVS9jwJQKGKwlJAYFZdEdhmz7ZV8mo7TgOeS4ohjIPrsdyya/O6lhaiPo+3VGeFL/lREv5kn2+0
28EUaDihe+77WMRrVqNQEU1PsNnADti/5ca0XQkxe6yFwsbWUKbxCUj7k+CA1YUXFt+xmxgbT34z
RhyeOv7in22XFeT+n7LdEzrwU2pnHYNTt8868HB1l8xwfzrCSNO+uc5YlnOjm4KjnjMPqK2r5i72
eg5DF1wwPYIxqXKupC84IKmTgBKlaFJQ8bTPe4vcoBJ34c+69/TxcpHpNfhqHUBpibohuH/mVEem
OxGXweoLkIy4SgUqd4tIJLv4bnVe0jql7pJojqzqartpwLsZtPZch/0l7hWFtk4NnMzmDkOTzYUG
IYwFlj+hgDX6+yIpDyaCUvo3N5nFjB4nryVrFA03c9hUURkMr7qNkRCXRnyDgRoiiFiWvF7gfcs1
XgARIZBNRsPYM9u8TsUye9VXIAd3BYpXBaoQOGe6EcUWwkoTaqyUSlAJ8k2kqs2uxopNeia+6wR/
a8sQoQnWZe4mFdivdttRKb11VyhvkNuRAmWY06+Zjdv6lkl3Rag6VlT6JVcOHrGLZiGAJ1Sb3GhK
X2hNuWGJpDYewQqLkN8bQT+QfQuGteoEUYGH/YT3L7NsGGW+yUzUVr4gdI3CldXk5WVmYJbMjmx1
ExIOzePzfLS1M+iJtwVgs89L5yg8OIr0WE7Bll1SSv1UoytRgH1H8bd4eVYHDZsPmZHRxFtrmHrH
JoKWa4TZMMhR63j1spw7AOHYb9Ei1/MCrX1fPNWq2rxTmqODaHMsQc9YxYP7Wggsk0yaFSiSBPqS
lfTPu1vmb8sTtB2eW+ElZSAxbhqgHK/Sr6KdFs+BvBFYVDPzTGt+gpuqDBqTjIQL9OVhH6oBxRoK
RxrNwfCSLJ3HlwuVa6fo6VdvTMcFsRKpF/RdMEfMbT/HdMfZQ+TB3VsA5Qa9aAOxYuEwUOo8cBta
vSEmB/bXoGbzh0w5D/HGPBDVmF84qfdNVBt50/owl1Xbb+ZKiI4z9HWvCq4YW0nsLP8gCL1M2moe
Npamx1jFOqtRqq9l7ig8OE7egjGziAP9e2Ij1WiT2HZbap3Hh40E2ZFxGaIi5QYkjsurXVIkA+Nx
EMw1mar2tmyWXoqH8U9w3eFhR7qa2UwFFOseERe+kEpeuWQt2EB9sC1oEziu76zUdnfG2Nacb2xg
BgOaj8oAB28lWgfkQck13jBE1/wker2R5xOSAagK+tUP+C3dz++Eb9n3d8WsMlIXatrDO5Ax+h7N
3VN7tXY1aqI9Yrz09MFMKrTKEC8i2C2nfK9fOvCoD49KFj7MaAKFsg3PzIE2Hpm5DCb620mYLYpS
9VGwYcOzSVsQw7u3VkyjWxOLUw7SRcJP8ERKoFJRmsml+Z6vlcE2GIxYffCyGnrmGyrpmP8ywN5k
jjReT3IU1fjSKRXzwdhZe9Na1euAjNbDG7VGMtEyTi+fsjBNBUlDMLP8PW1YhH2ZLq5uBpA/Ms+Y
MEkMSacHm50z1nHDhd7O4/zfUEHZnAq+/v0CQ6tlblDNWdiTddr6adtpm3jYnwbfBPno1WIRDmej
4Bt81oBh8zapmH8TlAo2VN7W+MHd7PCP1yBjkgg/cXmCFruLVTjBwbCmixqCsGthgbgMbEzw/BAL
K/Sm8YzHReBicN7rkk6J05vM/fJi03SuCXWF42MgvHw3Iy8B5ctFjrLPVqDy8Z9XX14ZrUVZq2x5
A7MBHeNJbeEEFy3H08RZOu7z2xIAd5cP9x7gENaffk6Sv93OBRGnH2ONGRfjwhfcGrZrZ8T5ukLN
r9aL4bzc1TV8Ykzm07w8gvsX9a03TmZBamt60gb/KHoJOFEMXgWHNIutLdpn0Gbm4M/bFAvA+0jW
uji+b6+sOQNhBHboyhM1bEg9a+7ygZM3T1g+8vpAWC2plmZ05AI8GcvhmYETAmAzIVDHMu3z+TnJ
L24nBWI3t0DwlxgVaxyssYqU90B+pNKruTIJltaFCw/AqDQ/4T0naEDkj7GakASoItuNOtd6/PvN
s+AVuEba1NW5rmrYo3v9+nMZ/XHggTmPkATBvVJPtU4Ca6TunPmmBpqFsqX3OxIrQtgSTkbIFiUt
igJEqyB3n4x+xBqC9835U1XH7NwkLZn79UoMik06IQ7S6xpmW05AUtNaPRD8lot6wDT88rgUrb3A
kk0jl8w2BRiUP23Nq9LK52+37Mw5KPsTaOKlQdbmjMZIbqaRdGpaVVUhZoIfcHweo3h2mr0p408P
5BjA6XugTVpy5JBmVPohkNx6qOE4wPoZROIQ3HRhDzePIeKmhhZC5CAiGwOzZ4+CYdYO9VmTS+SK
ColNjngOfrBScYBDHpr2Cx9mVft07kOJALrqMxuTdXut8Fc8t9DfSuLBWkytxwLbZ6BLAeh8C4Rh
3Ij1lC09lHpkCN2GzZbd9tBwaz6IgTbIxXB/EFQHIWISq+6x2U1xoAUuBHnzB9VRh+mKK5H8ynu7
aowQB+NjTe5E39s8Th8NFXk97z0U6EaedGTt34VJDDcjgJTdAj0thGi5PqBX+WGfsTaChlMi79RW
aTX5f5BV2s5dKpUaR25IrSy2HR9/7qOEB0epfR7AIdvXctajsMDz6BfBiNt8Lde1dekhjwD+gFmQ
YoaH92NET/ezsm/NTVxEio2+/N820uodXXT7ANpkvvV6z4mDGD7skRr2JJ+WP0ziFkdM4mF6q+7t
ll0MROTc1E7QWTVHSQKb9/OVCLfJAE1li6rh3jjKBv5302XE5DG+1o4Bmxjb38Oij+bOboBLUyxI
0Vb07Xs1b1H4UGmBmyb6hYletbR4Ktz3PP6BusyiA2tM9CfpVZSv4NEDFLmznT5kkb+eG9xe4L4S
gQohk72/alfPcpkLAbh8hZ5W7m+t7VjMA3DEzRSW2giHoyKOVu4ZI2rC6sNT+EMLAHWOiKkPxgS4
kwDJgdQ+fHaEdWN3NvZqOqpcUQjY6Pc/DZ8uYCLYV4emY+EvYcVnmOgf0fALLMlSFXT3FPN4DHuz
3ohCHHQVlNH/ovhmD7gu4bHh9DZWlZVs9M4lRwrV6vve8dNJWSLEew1Tf9aHcEKFctonCy5f8wPx
fOhN6Db1W5WkfKTJh8FVkQyHd/zSwZN/drpQdCcFXSUNqkJQ8VSeJFzW+h+jayht12jJIJB+WJ8u
cUWLci+gQbdG+z8KGag1DquD8HcF7f3OMSiwAAG6vRPy0T2kAqxBKyD+Vf6HVpVDAawnxMI4kemT
aFIwfNoeaTYzJzWpyz5gl3QqYVVYRH3HGslXxK7/KOp3uBmWSJs5PzSwcM0MmW2iKy9AxWf3vIV4
6KM5xtTHBNyRG9fEJwUlfGnfCZv/yL28TNCD3DUo+LorZkoTiJ7wYN8gzvOGBxhjuqplAT+v1u0x
1RZSCEUs7LCd+30VIl2MBg92KyosCQhMuiFFSpAcGuYmHaS9WxvhnhCaGMPODsxXe1yQtN5orjjf
TVmhCIbZgauVB/EZioG4lwyI0HGqDSasljY28v5L9voRDDBg/vmSCU5VGVnRQtFiHkjxTcJcSwKc
ZgNy2avMcRmE+eClgxJM893XDWDVbmoitennGY205S29LbuXP28sl5hfhbSSBj9ma5PEY0+An4YS
9WdELsmbW0v4LM5cuUJysJPg+Z4XZtDvFpxVcZeTav16BijSupxldsoi4luinjeJ5AIa6ZeT0zp9
IQlNCFc+dgQ+zUm9+d5yLo1zz+r7E/yuKVHLHTytcK9VghotBOtwuzPDkq8BpTnAINBODww9+7IY
Sipw7fxnnGZLmu8GLPNLdDe4HyyaAva/YhA7OCkjejtvu1cv45ko+aaqzJv+BQDLw+qNkhsxLkV3
82KQXqbnso6F0Zv3vX/ubj5q1lrsMY3XCCPiyMGVQ922X0lbILZYKZidYAqNZ+NUo7YWwM14S4jG
Y3GXJYC2ySs5wE4Dy9nGzRzG2npjzFtAVwDvRf2sJJF7LYYU2lnZX/T4EZ0H7gN5Bm6Tr3KM4iGQ
8Xr33U3JGnaHNkMjGm/rtOYaDFDWuRQO+kS/rlEzG98Un4SoKtDnEa9DTELxkapUEAIpWTdFCtSj
v4R0fjTy5Xy0+UO6knE4k3/QyHHyBNH7y2CRIvB3dA5/SGPNI12GvuGcV8rLoEJL7LgNnAwrDkuz
hAepgviaYJYpjDSKHK1P2i0orxrv1aGqeIpbhtUDKx7z9shw78qD/bA4+a4b7hMH5tzVeZGyOp7g
me1uvYaz+v+wnlCbytdFTuz/gcLy/vSQ9650d9pzdCDSEcZkuQ4iw78fhQu70OS8dQ9KWA4pzDn9
ewe/pPhFgTVMl65HbltpeReoGEFnHqcT2EDjuv3GsYAW9dg6//noZz+/+wvjzsujt90b6AQPOp3V
U12u6uV/8+vtU/gdxbRn17PnGYBNT34Z9VKrZkeaGM7gzXLUvX5q0yXqAPpmRvHQP+D7JqGxKwLW
QepI/VffR+Q9hQwjud1o+ixHf31q/aNwhut0b9sEI4mLTt8QY6pn2HtLR0p2x/l3oV+SByNl1q8s
5uwAPQ7E98i8llrTVtnul6xK/BjMxfFa1+7ihxrxL+n1hIH9EUWoWwN7gyaWSkfjXUZxM8Zvuyo2
ULtblGkDCIr7idVBC1rVP+lAg9DRCmfAlXwwsk05u0CLzblMmS5Z4oEEgX/bpXhkvP8vZKZVp4yp
jjDPijGYjNNI3sMQOtrmAv/67wINrm52cUrhnV6DnGzRD8meWL+ZpHZmR4cUOzU1roTSFfJP+iyc
wjtUk0i5qcOLqkC+UTbYQLXssnHKU41lNRu3KAvYQcarZW5nLOzArMGKSWdl50g4Pe8oJtxkDGVA
UuYVeZwCtm2zW5QGuiF5JVD6F6vtbNOYB+LfoUsNAClw6wRq1IYJpFF3x6GJl0pJhgmdXtJAesIV
tHW1aafOtocyfvf09Xv+US7ZGoQlwdlRwDEU3DS1Vzb/cw9DGm/lLfM3/cfH2qrOUExWNeqAP/Qc
mbITbypCGrnS72BYusdpg5TNnEBFLESn6Lr5e66up/qXo9iomQ+me41EZLBQLeeGBwGh/QiL+pH3
+O1UIhrHjnoh6dwUhlhHZA9ukhnidPqCQHCVvjNjjphDUqfFlWzFvraXbi4RQaAJqAN6iH780Oxf
4evDA8do8yFixNC1wsErZZ/QRv5x4M3+Adja7wAgMSz/Q+W7NUcyvEBPT6ERdMhaOViXBx1z390C
z0CYS0kgvymHo89jSf73EXdVoqaTRfFvZUCnGg6PW+TYmxSYzGEwnwr0w5ZnsK/mUt/TObHI7cMI
44v2opDldYHGi+6inXdoJKSdMiImwu8B1zdablPr9Cheko2DAb9+8hLRQ7UEcscIXn6yXgZiqoIB
ggOXzN8lFulTMP2Mh4SzzR3Luw78Ccbxafq9y/sEmP/NAPUIXu+tqbWV1HLf6ZvmPfmx6nYwV+fW
Yim4ZRGyUkDa5fpiVQxo32WK+QnpMhOuS1JeP774eSKzHCFXzEV5UhUI6Qj7B4aZuZ5s1HpT03JX
lB5ox4qZXAzmstV8a0VuExg8vXWMRgOSXpmPOyM4S8GYqLQkLKN+HtPUA7MEZGnXJHiKnABDN4MY
+3SoGNR6AQDWaZpJZcyBplQLzP5/KqndTaiIWT2sQI0SbN1lifn1bkR3j9lPUbgyyy4RBnHUx8On
+jBSKv5dQBhFYOeZV0Mo+V80ZX2KE1F33D/gb2USULlSAtMTgkti25/QpiU1cg6O/4Yfr/Q31qCB
52F4BnU95CNpF1/KI9oavK0PWpq7FBKUFh5hpIJlc6Q6aaH8XsLpquCHdCApXPiJ1bZDs3ykxssq
m/06c+ncQhHp37iI+Aap3GGTWyZ84M9Ll13Vb7h0LriDf1IoahLkI4kkJgaij9acK/uHwd+C0L2R
KB8YUX8wN46fggkOOTSY7s8qXLxdTXztJFLvLnHuEZSLZAX0kdYeadP55QXvvopzGq23IU2rvhjm
x+YAK6VbszsIe63QhveDpDTfyPwpWuuHZWXJcG7Jw5ZJtjoMNVvih8Cm4va8clVvDvH+6tULe+vf
V2Po05+Lt2Q6Ko8l9gHoeM8wNY0I3eAFYd4uKOwaBBZpa9g98jnDfn6uxOlhDuI83mzuMesOh2cV
8xqTFJz7om+OX5utTW/kdpujX/wHRGmnlHntZDZJSkUHBF9wAntgouleVCdYsjN9TZr1ByRbeRPy
Q1dLF7SlI1ZEWw0J7j5mO3sb3C9CXw0XPErpwGXK2HGKU2DyOY+HVw2TNjuPH55rsnoAzvUtUM43
on6gmSoS9EczMFq6Nx5bAAvV8NVpme1Wp/Wul91R2TsnSbcOvE57KnhxNt9DYAqS9N6tvRlGii6w
dhaIq/B3JHKA2pXcuZdcjqtfRZNS2SAeOI5TPD6QX0woIS93c6qMhurL8rKWx7M3w+gjY+Euotyi
YIQsewvPzz/9jOFSltuSLshKcX98FxoVg0pu6laeM26CAcm8ynXut0esHV7KkbCVowtFDthltZyp
XdYClIr3TjYTMVRovzOI2mDosUMVMHVH4lb2rr4crPFAGPxpwhLABy94zCpruzOHnxDzVT5XaYTj
IFY/SvcLbwxdeMXk4JEuSyTb7mDG7lMQfXuSEM3bzGk22s2qUf4wegaNvF0AdFx+UWMb07S/XV7s
ukJ01t7ca34lDBOEd+TV1UZ36npf5bisw7dYfcLJxmRSJKlM4aBdaIZhAP/XbDyO73B0oYx/6uPF
KOzd9YDTANlHWusPSjBijnFOKj0SQHmaXZALSNNlN4la7skVTS0517xyG7qmfTuii0UkEyKT6gPX
kBBMAWBCR+DGi1RwCAu8T8dVvl/8I1S9mFN6A0CF6BUmMk1sA1niQSmcir6IaRz6LDBHt8WxqGaL
JC7FXr1Mr8ksA9XaYADUI/7cw5H7D+ToJyhrAomyp8VywBDp4SCC/CBhKhxggOJOpVdl4nTpz5Kw
1WGezLLi6K5ZUcmI7dn+u76EZee8IeNpGt6zakQHSYIO1GmpVtQccqIQORthhtJ8Oo2r0xzoKwVo
113d+ofR6fmHSlC8VF8GwWYr9qfNpnakYVHDHVGKWsye9Bo+mEKmP5QHIgWkLFQSdBX4wOON/FFh
p2uqGbC5G+GKfTYfGrIlbxBXWxAdwVJwiPvpur0+ymS7WSP2zMk/Gvm0ckShtz1qroNFaQSQgZH0
rV4HYTMAS55RuMNdR79RBwMSsutPOdxI/h7BpgvP5FHEV7/mIBCaSfJ8v4oi+uYGi8jWJYrGf61l
VnMTz10nHA9VmwwC4BoMPyZ+BWghag1odilXGjKb2afXcsfjOrwJIiAlmT898IeK7Bci/zNta/jK
zUTDBUZJp8gfxMhBXXWz/yq/WRQfjV18O0UOBPltFZIjPfCVeRRJJAe9961BrgZ2vtCpEuEMt8+C
Z+ltImDACylkklRe9S6TOVxQf0VF+nxK141phasqdXr9UsZ17GlY8m/SRUdzlRc/Yun3x5gP/GEg
Rb44XVzZOm6vdIT10gtb7c04VvF1iZzRFeDBq1TbSwq1RBXSK+gMBbt45c5FyjhGkeUxkViWO5TJ
8NOWtJde6VXK7BOMfXUpWhs3kEk9VnI//IBecVQUDcfRTxoM2DtAG5B5fcFLRhCcgIr+c5/wOo4M
u6IOlVcvzIDBVtAvPOf9jr3rlc+MRvqUs/kDTp9YfGcn/T/oY6wwhYPEMt0vX1RBJldzFr9krn/5
zLICjK0bdD98orAgLslOtAZep2e2yzETh/OoxhPMp28nT1FZBLFKtuIPrikzwClqBI71XUcYhhrX
mFI8IYKlH+p+5Bh2Q8Ilrpnp7DLDfnzMgCmzQoCSldYcAJO0V7g6yOgOfUTYM3IhwZLjz6tr1CGy
5jFkGcVYHFr1158fE0BgsHGiwgWp7yIp5SAI0a+vdBerQ4ZaNPm2XLxs4+2JXnvr6HyG8C6bOba2
wVcFyviiDJxueMgLHAdHt6/04Dbnd/qETk+227sARhwJzSsf/IcRLg/VEhFtdlr1vquxB8edAH3F
DRyMDELW54cpRpiU33PkfcHkLJxrHzvOjcnk6WE4F7wc3M86OXlybdZuqLe7rIDcFWdZPCkMBSeW
MBt8Gl8RATq3zcm6dftyKoZ3iTMCsSzcvw9xI0JEr63l1dBqfI+UQ5F0Vb43bhaTsfRCunZcqcfx
uYEI0ur90gRU24Pz0dgyeqTdd//Fve2g6LRcZyPCPWEGWph1OZQd2vsaCd4FERf/ll/sONknHL8m
FzpJ2hpPxLytHVZ8OvD0LL7wxxJsouTOHGUoKZf+5jZ8YBxQUw+cbMY8KFLWz0hihzXyM7XLFsIi
BcU78YZ19TyAZSCKiLZz6Vwq0qdUyFjLucQufZRLsRf9OQj8BHsmc0wT7bgeVSbwHxwIYStTLoAQ
GEGTnkCM6MV9cHfDpPsdQV5CLFiyNnvtfSznPm3LaOCqXBO1d3n3LXISjROmWhVULUjAMmIH4WuT
gKhWZPubkFan3vRta05IDdOIy4/Ve4MvzMqHnZDzpWc4lbVlLRcIQC8cAZRt3dAgqFOW+y+yg60p
bxInR1tmB6k5PaVQHIE76/gVC1ukIiovAFYNM8RZQp8tvCJTf/nj3ZAXo6RPMi0TIw0tBYgnh1dE
Yaoc8p2KZ3YuADfGNC2NqC6L2aBFTPqqoSCSbRdhq9t1kOdEXW9gnuo+WtTj7eBUw/5Ktx0ryvfJ
KhfHli9MkjISOR5YH2sdT+sM2WFp6pbtnk/EmzcXlcnrJoII7JkqcYnBErH9+AK2YiXmYrbrhzXd
eWewIAAYY4Wcgur547qkmuHVx5D0o4kTy3/JVSnG4Xi8x++9GmqZJSbTb/oVjxjcRG3oOxY0ZGkW
xsaVxCZl6xWWEtIoo6ePCh3KdPkt2+d//P1cAETBkguZ4yjqmScwNquz/zpxdhVGg/cWkssyhfHb
jq0h536rsAiVfhAzEerETlkXU3ArPeLcEO3p4copfMFTUKAuDiuRzU2acybsbDlU7JgoygvR9y5y
F7KD37skk7L1qrp6Dw+v7z+kRv8zez5rpibgmI2x1nrBLSPbDu97NmN89FyHBZcv0NeintHhhlnd
dgJjoAEEW5AntsrjPXxM9zo+wp6ABXJQhrSCb8D+YUvO/OljO+7mBiK4KWyw5Ef16q0GNBjakQ7r
3Ex2MIGbrt522wiKJ664CRe2DIJfml9zSYSeXip5SPXZnC1KotGNzF02XnWjKNBTTrbOtoF7uLpY
21/FPZsQozz6VMaqZeSmqcMBZhTn4+fJkh3Ay8Ir9btobRZVe+XRhr1q4M/Eai8ioLSpuvODsPd1
ptyxut4Oc3A4maLjubpz739YhvOJdaXAhgMHNJhxn0VRwY5wsgxLYIHcHbHce7vMy/4/pw/NRwGp
YZgteEGTqeDukGiLkhnHxjiCWRZ8ky55QxSlOzrAlmZTu86v87ErZ5z8jzHYmffyupA1O5Ni4s09
ezYq3iGiiAjXDHCcST3fEup6bArTnrkMyh4usOk9nd/bMtd1JuuYmFKYyHQkOpy8tGW283l8FsJk
anBAIwFProScAfqnAO4+3bgoEi/+pLkzb/Gd7DyadATOnqvP+zQuiGbJgnabJ96HFSotI+QnUR6Q
LXvupzW9iVJixiP5+pjqHHBJE1wvD2KYinkfNajYxewK9NMF3iSAN5OeByJoMKIlIdRQw+Cr9s/E
2VyWuvKgbx28pXrIGq11OAs4fF51/RUrorRf/GGfOY8wgDH2nu66UNc8TsROfdAB8vWOnKJ+1yDV
a5bWTYyvUNVeAPU4c63OzJE9Dx91y1B2Pazu2R3mUq+yYnNnyMxVCZK1Ug/XLLK/3xLmU6xgHocV
W/A9rBeEfmJaBky/8DPhf6azdMRdBknThwIcB4kswBzY03+HXxWNkypldkE0SiN/hfJtStMeeZHA
Cq58zmGSVzKcbI+zgj7AWLxUF0JYgA9lrhXRhPYTJ3mWeWz+Bti/9Z06jZAEemmo17r0PKIOTkaw
IiAgzTXCkjmrim+grfoA2CxEwAhCUjIOXjqFsAQbMn4wb7NIZsS7V4INq3+TmYA6aHVI+1grTyzV
O01NMBy7Cc3RMZwXPciNyY9n4WOGj1vele7fp9BQWhiWEbB1KIK00/DvTNcQlInzFy4F3pntr159
DPkkLLgikJMTh5wqXDc9KacuybLEdYqLdB2oVnVYLtkPF+U+TZ+f69eXng/fanFZ3tgEhYzRACeZ
5lYCZqrajsjuowAQINz3yg/3S8c/hPytpns5FY7VZU66dmvlj1AuW1ywBIpmBQw8SBKACFgMNx48
5BvXXLlOPa5W6K5zVCvXLu0oYT+rsHQ6NsRs1qjXM3KjUVOpl84ZziAO+oj6PhydYOSur4OKREol
pM6Bx/FcwEXN2nsPFdUYQb8o5SI6sMZHoSxTARFRs/2DoPv4UeB7u4Y6TFBoGCa04fV4sKIDne7W
9z1klm4iFAQRBOfRHUxSkhF+aXrW2CSOhGf9Tc0CW5cOJj1jjt2u9tdxXTip+Ase11yGpgOhIs2Q
7ylnK/igT4tt4mKt2vWXZIHjhnz6CPcm8yCDt6/uT8K2fAQfRu37uRpKmA0X7Mf7iFJsV6Bfd9W7
Qy/W1B4CpXtMT/vRpVGSd9m72eYxEPtSncYYaAAV2lLdpaywN5k0PRD5MU6pPu892dgyNXtXuVXN
lNQrkk2CBUDWTV9I82/dOKCJujTL88/y/2eYLh1WAZVkEwrEEMcCgK611pBYzaSFzPCr87R9z3it
Bd12C5FPU+DHowpHlWcaEwIpWtoAD6VlgDpGLqTlnW/20DWRfTcu6sCyIwK6Bd9lVS5G8AjfA/o9
xtp0H3q2R3SVVxTyk4nfx1RDiAtCnK2tR3Ng+8Sa7y7lQw8FBNDTQ5fjN+yYwTJC/2eKTRl6y2BA
6gkX3WGR/4U9pqH6crc44lws1VvXRyMbeKu385KDZ3qjt484MlIjut9NT4sR5d9hcif1zhby4x44
5nIJozYdZDpl5/+cpECuAYb2FoE3sC4YK9F3BFakD7Yp/narmO45zhRpa95rySde0i9EI3MUOcJe
C6It0bzqwgsCeODWijKzIQdM2pXozNOnv3GPfwYdEXEEYbskukjO/oKPs/hUhzUSTTDPPtFnnRK0
cevPXjDWDiVOKNPxZS94V1tO/bcxBSJKSnwgK7LQX/VDsOqbvkx+QhZfMkC6p/x881iUoDYyOMf8
5iPGZXoSZUu2O7GeGK/Fv8KS3L5i0L5YZ5wM8OvnIBmZehZ+7YyOapulDv9aGCrP1vksi67URVtq
qtV3EjdKKinnHGOj/ZMB4Eo/4iz/B6Bz8ePm3aOEfZvTwuuU5BS89y798XQYpyD8LW1AS/CmOj+f
gNpwX1TMMvFh58mD7hBs/8fdJvRXZ0hyLaJpyOrXn2YhcDC3XqF0SRAV8y1ZREHnWzzFd0Atqy9o
mOJ085SB2JMY72mlQbfI9uO59jSAWl6h+rRfFXqrqIZPSNybfG9KYvLKDN9FGroGXGJsOJ2TNpvc
6yiT0bYIdJdjZEb9X+r18pNLPzuOQj3OzMEpTKP/rNNn3mI29he3OpBhz6Cj9nZ2it2GdD2mKdno
hs2BeLG0XoJWXMyY1DNDEAT7+g3sxN72zciqw6aMz6enfbScZAMR2E5hgaoC9H8i3Az7zpnO59Yy
3HPbhIadryQf3yWdNBztUbS3vg1tlSM680FfR0jHk0qVGjNmaq5tJ6V7iABJe7fuDzXznnwqNXv/
4ux8BSYDhA4uC1O7MUPlbdSVjAE+iVo3hLwRfmx1l6MCQHjya4gmkMqZOdNbjfhhyrG33yxawnj2
1XsZ4WcfZX97jB8vt2KvAN/6ZFjdiZ+vEUWNnScca+wQ0mrmvMfTlA61nC1X85R7F41LrHM3bC2v
0BcX33ieJuzqs5+ROGgrHi7hlMcQIrm+yBKcAfkpa5kSLRnP5KTE/cOsZnCBXvEggP6J5XzzinBc
bt4DUYjDdEG03NSLYDuTiV7HHxSLRnuSSthTg20dfmpwiMU5PdhxIo5zoDF/QGycv91lw/ESZRao
tCsIK6I7KViPQKQFA/4SEM5IC1Lm/Acb6n+4ZTbpwfxpb7gyznNQ8k6zVEW6h0HxT/A54+MwTy8N
No9XQlbWX+YZW3yHba0+QzcFzf9nXG0YzIvQtOlHSxeMD25PenIY5XBlZN0EkeOWpjO5hVV1wNMt
R2Ogab1RTzwWrwwky0EqDPOsnhUZ60ZpnT/2zwvZBET+SQTplfvFnuLS4HnW/iE7KgOqmLenv74S
PuV626K7uVWNJPXbZS+8OnFYueAG73R9cld3BwkFj5FBy42UzNCCJqGVHgorHOME1i7PRJa4hYi2
xGyXus4LgVc87lyCY2SMsNlmdbi1+dXfDS24QPw1ja/SdXYRCyO1yH2AESb3pLXCPj+WD9vDmTab
bafEwAcqs6eowZ9wLmX1JRFK1odZjY6ty0JDnpfRYJP+JJ3hfVlBNAiRxVUCi4o3SxGfsLjddsrP
XI16gmm0I9qE5pcVo8eSEyNDhn1NlrThS22qVngIIT4CoZW6d1U+6qAQzxuI99SxJxFvA9WszJoZ
ifcXqi4oPgoTp3QI191sKqC0BDF15qLR8iUSy/2URxn/dMui/uIqeekK4QYqVmguCDQztYYTrwLF
d+JdLlg0xV6BRQc6m4Aaki3NGYfjMsQO218+cmU+3a79J6LpRr9aryy9qatc45MLV7rZlzZy5Kdu
0/0gKxYr2EuIS1PanyI171BoFNYIcsUBVbSRua/KL2nuRQB42FuvgZzomB8PKdyx4kaGdh4L5ikE
HyZeY0NXhkKzpxilikG846CCc5gdwW2iFY2fVAQDXo4eEbRq6XJtFxPXfpn3vr06bBcJzB6UUDeJ
6BDEn3k/Ngfum+T1dxNXR1ocEzxthyLVrdM07EXk6DF6YNPSd+Bqkce0thFBHVctGAx3ImrOdtzN
G7kNSEtyJcAct2fYvP5aWrLf08Na708XgwFf7Q6ZmXexEJ+8NWbyTwOMvNa8s9pkEcTVJyjOd4CY
B/VdylP0e2d+8Y+lm0+3l9HfhGSZ/7orrn1NfEJ1E8vstd+35CBU6SgO4/ha7GEoKgSTsvgtcHvf
5gaKjIRVjazmQ7BrqEuwTshX8121RS+i6E3OufvJ0v4YCyENUNdCvmdJ3fDGvhTt2yHlNApo2xx1
/zmnkpnARYI79LCWrxuQmwM+p//lgeKhY8ToVtkt1bIP5W/ao8W+psrSQVv99AwURqAkfFfUksoc
vSCcwE6LYeUirwdB8wXNe4n2ycqbrG7dtC4GKA1Dh2kAWQaL9HkJf2t9j2YUW9GvH2iSncnhXR+5
UxNrQavjB80XIbnGMkeFXA503F8b8iD2/5UvsNnee2FXQJvGWPyELkW7wISfCeDg74jO+1ws/wSX
buqt1oPzWnA7o9/r/KDQoJU2qLoOTmEFqkU0Q2iRbDmEQRYFsgsE9akfA8uWKVFmc8LedtCV8FBd
D0wdkVIPac6YF2FZJ3PTR2MlizEfactWY2TLPWhe19DFsPYVHZKxJ9O8eHnCuEUBVfaTiO59seW0
0iJPwSj7WZ5t2j4+C6KLzkKmatbcexy7StI1HvLpJlt8VFo6XxIc2tcHgM7OJS69HSXb5n33uEks
0uRtBM+Tc+Z4jZ5mVbpKHNlV5S389cuVvNCmpMEv0s+ORzfUfbst9CGY/cU4ldKHb8PZt6JaWChD
er1dx2F5Y41ov3I8NseNokot70lsiIpEbxrmVPvLzb6bHscZRqvNDknk1bPheuBHh7jLYyxMgEKh
yhkczK64uCljRJYgMxnIo78cfVvndsBUWpE50GtHmqaBD6ygBJlc/zCQL1HZqJkNziX1uWBYcHQB
3WzMznDMa1m+oNVnbTtDJvaGFZd8QcY1ovv2U9RClcRLX2+VQxSyDD/5XbVPQHneoH20kT/WzsA4
M6exLWNYWmCehCk7TKrSygu6IR+Aelv6P2zr4juTA7GwWjRrARMZrpzddFDyUx8rUr2nXd1f4s35
+lN/j2yWgaVjOp99QTuA6a/SqUOY76NCvItsqf3yEdXJ+0eLd1vIvyKGWpgIiiNaoap5GTRZHHEs
IATI9WNRM397TRZbf0rUl0uJ8a3Xu6yzInA7FWvRn2hm4wwuQB3GLZYDevhT0y/dZSbJVnz1mhlD
NHUQI5m3Zb3JQ9gUalXMfwL7qnwm/gWehFG8Os7BFiYoZrwj51rXAb+JFQwy3PUdTFX/ZMt+mTny
VOUT8YMqTPjNoUu2VMFOoQu4p2E9qByG4SOF16GkQkMYVyca6OOzOSmuIpkhCMWtqTtH5l9sKItL
pccZkdlYUr+h105qG/M+xQlgTKjRqWzWpDcLxrZxy06Tsh55JZG7nnRQX/BEs9PQ9xMCjt7Lgh69
fD0veBvAZza585iIn/ES0rM64zUzcBJGdksDsYiYHa9sbhZbpmfRJMGyqCH6EQL7I5+VQ9k6RI63
WUSUa5/DdPD40awo9ZfnGRh6UftQ88qIc/XGfy4JzK3MR1/q9ZcYshJsiXVswUQi5SQD7AUvNRzc
hf9a2L94CbuiTLO1OzQYwC0huBRse+Z1JabY1QkyV64oeJ/rwmhrFguyOYLgBmafWNOr2erXiaTl
IFtfixOAMYULb5rrtvyBIc9Ro8Y+X9ktW/BEJvWglCj820VOTgoCZGa/Mz8m5bfh46BGtl4NMUM9
uOApLPAm3KmGGmVG3l91iEdblkq6XHy6D6vNlGt5Ab4MdCzxrBBPbJbEd9UAwPL8Xfz4NufVJPBv
S7L2xahxBDlT/cgeBzajxod6T7t20hpii/V3YOKZerrivRAtoXV2qqaxm7uXK5dolkLt8MLSAWgb
UnZvYg3+ZkA/BJ3nMcv6hkseBa0Ru632O8zMa1fM4dgaEok93wE60oKsIBEB3RTM7NK807h2bITE
nhNYsTbifOs/4bxYUDaHJzHSmOQPiDVsp4cc6Mp5HvFcxA/iKcOb5akKjIHHD2dLGh9T7LoTsIVF
3QVCTR8xlgxT1k4hh25NXv2rOZo502HlW5IPrSXPRJKIInuYTdksSYg3Vw/6btIJqkN5X39TYYmF
HiV49XwVzD1g0aG+X8BOJoBk/i+47vbdiUyRso0OaP2URoQ7o9E8QRJXpZ85A98bZbpPstfMTi6s
3gTMyvJeue6G2Cb1E9WoMT6r6OROXdDZW+mgQJUCaLG0JzPYEHXVhOnMilaBX+ynaPl1B60vKj/F
6LhSeQJeVbJq7b4fycWoV7t27FLFhiMkQDKJaDW6L/JnpvcdGgQ4jmpA8QO9w/WEEpsvVUYuyHFA
1EK0ktnpkyjcC2nzz2572+X7iSw8oqsFzXos9tji+UkdqFmk8O7983YZM85S+nWpVa22f36cwojM
+zdX1LTK2YxHe6Mg/30If6oPb1xJMrGOSi6hOf7o4NgmyRPwoXiRrMJaonR5pw9o7EfWP6uQqjsN
njNAJ5Qp7Y4Lg2W6wgM9Wr+cP2XSTP5bdZHdRmi00jdmGqXA4iHH79Esh5z8pzfyR9E6YQqHjf2T
z7LZMGslPWohfh/zpI0cxZS+N/O7gDCZC0qQ7IaB3sS1FLQU+d54OZKF3stKC0WzkOR+/3ouok3k
cFdvY/GQRprNEXXWSeym3cFnpW6zmqpgoposcJqwQr0oBBipwB3ZrOed2LtK9cfLoFJWGwZqUhzs
Z9byYgDzd1i1wEzfN4gHcm2vyoC3PnJlK8QHB/IsB582Q7TWKC/56tsqyDCHvURkP5/ZWmXp1cnj
ObLYSvzbzUWfia1wS1dyYSjnsl5Hs93ZX1DodvwEiCRtUVkTUj6JccGcUPd2uFocetsDBqlvsk01
vhM3r44w/m4E410BCqzUOMOPv01bAmqnrShuu9HLpOhvkAMjcMqmoIHBozivu0qeyEloFYzsRigh
fPpFU8GaOcH31ddLxilv5YJM9kuB6oqvdeteINq4AAy8UMnuXQ5Klu2S9aon1imG1spsR4rqmLnu
liUynDTqc1ixRFmiEPjwle2stw3x/47SrkHoW5nAPq/e9ktiZ68+SCxMvbY5WGx+eBRxenZs9oqj
kuZYHfomoOrtmdH+Zirhn507o9HURPH95gfNsLuK9+phewZa11T6vQ1iTVx/NmTHVZF7rrMTaDzf
/3/+BQIde+az5RSEuynD7BWE81eHdb7NVKTNzjaL9zewTmbhw3Is4FuWzFmvbQWfPPPrzcB3ChDy
QotU+ia09Pp0+ZyFFgYonvK6f4qNXYENW9ZZyJvbpkfK9E+9Dje2xtPN7ck2ZBggZNi7gZE3CWSq
v/tQQf080RcEoqjaD8z+7oYjCLEKRDpD9OGuKjogAmFg5OwxgeVYHehVyajAIH8b9447mvbhxrSO
h2HGEbgny2DNIt2F8E0N1kTRKeqZ80WmSH0EHJY6usvm4YsLKBD5t/pVwz2Lsvn2odRVeEQpXXti
19tc3zw6rCqQ29qPieP+n78PrzE8iFXCLiJF04npYGDiA9v3iwSr2nNW9PKyz7AMt6vTfyAfathn
QtJPURa+HMTYZ/jbDzEfoFh8NQSYhMc2aN/gKdieX4YatbmZrGsUMSlziHf6M0+vXVqrqYTZuCQx
dT3UmRIeU+hgcJt8HKIp11Vl6QYFnDtlgN7TwbqJ4y5P8Fn6Nd+hExTuP9hl4unBS21D91mDNFpD
Fev13sduOlbalvqgQrAPU/IbVbtTWAyHGgykPVZmafkklkUIpgtXCDV9T+Jo37+cm9oJwsy/IAA5
KNqaxATjU4hSKcpVXtKseHQLE3hO1r4WmOeJgYggmvCXeE1qmNwAUkAGPbg6d/J+8tCMldxH3G3Y
GdiEE8yeeA0Ue8Nz/ZiITN6TuiqX1SHshYeRwvTchsGyPpuOYjQTaM0fkz/1bcpQ4I7uf6VA1hP8
ymdIqWaLSrW5MLGnpzzVzCyBoMl2zkP6SeqUzmypYU/TvO9Uh0f7ZiAjbm71UFUAQL1qkrvuwiaH
L/GW44ngLHDG9KKHYUXoFiD1bqjnLYitoZyQELgxB0QETKRTCbRjwYl7TIkR9gSx2pIpNTvQGNBx
QVK2FWqzgbPQhqZaNLlL+1AeT0AkwEanXUn6CIEOaHOIHQViFDi2ercz+i4ENZwuFF3d6ycXGQR5
6OmYO9nynCvz8IRniV7UP9c7OWgG2xNfSdmXpTeNcf7UTgTcUdKIr4P8xnnX5nrknIg+3vD3Tjqd
S8M/tvseD8le+hgxjp9lP2U3KEw+u+03U8owCDpPwNasxtFRO2uN62kmi8v003Z0+oidJzQfNEZI
sLbNmySjPVF2lrH2lEWrdiItYbkJt0czvqrLQsZAKxQOpbcT74NPgRPorBf6BqvZKWoQwVCkRQsw
jrQRs2yJFpcY4i7y21t78esPLNP1BNacJboJhntCOuxJpFGJHQesQQw3jegcXY6XZ6ZJL5QMmblT
IuyGgWzIiZy4Ietf89T2K+JsuGDS6WsTAZMRhXvH2eoqMPQoAFbGma1XvlW2RQsuRMryTjY8inXi
mR0wzb1uBa49Ii39WkobCs3fxZ4ONd5X13bHMeC8G8QyFdfwx85g6TaTxidN8MQep1FDOKjCHuLF
+T8h9MPl4VIX1IFEmKzx4Sr3yScPkd9sqZMTcbzj2oDxszIXEFjNtN0qgsMzQy5Gm1Ud3gPRsqcH
FGZz3CMTaeHtFz0YldzGM4I0am/fbYggcVOUuKPEvsv7HenHiuJPVkFRE4n2WjFUmD/d2/Ijo4zj
J1MmZHfxuJAUDwMk37r3nqBGSnS3Hbut3oYPmJ6ujUfMTx3kagFR03vNfprQB6DY4SyMAdqNL9DL
wZEedbFyjnKP4etQW0Beq5h1FZ7nLdIakxVHe31xHq8GaYk/Z31vMTeB2iaXibJK1YCSgoq+0XZt
1sajGPJtMYVIuQO9FA+rsyvfPi7VWnk8mi2EmD4Uwf03CtrU8Bql06+CwrA/zs5qroekNc+dnZQY
YPdyxTQ0I2VvPVjlLJL8HflSc+sW0vsbZ9hmCsTexArb1Rk6nyEAv/mI3rqBgRChDeQKs1A/IO1f
04gwectB8bAY0LooYLnNqyr855hnyqQa/+Li3wv3TmsTR4e12ryH13Nw9R3boz9wU6rBl/tkH4Kl
GU5nimQIIvoLWV1/BrwEraOj4VJsh966Gn8sSdYhP9ofBeM4abRyk6fhP3BYHCtcAtU9jbcotiMt
hIxmK7j5VJA44uRiiprIZ6GJfycl73BBwglMFKGHJPVteS7qxdhVgkLvXbKf4A1Z/7orN6shxWFP
To/up6Sz8h6E5pKvJeddMtNqsRhH1aaS0k2tnQnkks5yDhbozWQIY2Uiuh0cEKooG1wKm4oLGIhq
pYlSeK1x6BU04pL2GFsquOeLn1N3QYymje8fah6rjAkXMuIs+1QYgyNRE6CT6QkrS73pD2e8D7vf
zD1asoHn3Ly7mx5bG0d7S9xgmIsLPQEoRw6W9bZUAZCMmYC+bYACeMmZ71dSnx7bphcnaMjekRA+
Mg21TvZsOT3vWKmap4uB8ZgPm/XN82oyQ5en5RrqE5U7iHQlXkqvgykK5XbfRfcreaVeWBU4IqL+
AGyqXOd+lT5nPAJBeSMNJhwZgJZLAjN/pzPvTeRZPAF35um+M9uV7NP2L1dr677RmvMcR+RCPsoz
cZBrS8dTdxwnEBfWdZsAfL8EJyqAKOSU/pykgdE2Ge2DxwUnNSSIHtc83ns3aZYWhwKhgG3eo5Kb
A6Fn+I7GG39Bof9cBgrIw8vaChlEPHigqb2YJYkSG7NjX+eclVv+pnWRmXG2t7XRserkEfpvwNXH
viLmwdBkAmGtATpT8DR1Fr1dy6CAVQyNvf4EirxWsJ84tbkG4UyXD4ljx1zRjbpFmYwCH24zI1TD
bZuNx+FvQKu1Qu9EohRWuNxhLRHIq4uAwF7iRNLf03Ru0gv3U6xPcaJAspa3HKiY3lRkoguO7UUZ
/pDeilwoD9sKQGaEGmsBAx/9rSFppjBQz03PlY8Gad09ABngwcOpePffxHYCrGyZuMRCa7f8jPc8
CXa0SjwrVepLH/1aMKOx6Mj6HUCWis4bz8bE1uTEQkY6J65gDzt0x/YBUjaz8CCYQpF6K7H28UE5
6Pii+GxKiuahoMi9QQW++UDlGMxfYwqE1IPeftF+GubVkv62sCYL04LUkj8+Yj+9eQ3wxCPHbQTH
/n5eUno6tRJCooD4keqd1ArQW9bnTCj/isnGBtT8mfDuMKsnrtLltlEeyP/y1J/66xhvSVVcbjv2
m7Dg0+N/J/u+5ytFnMZQ+/3xX29OpSgoU68BzEr5eq7rUpprtyuSE4kZ8abv4yF8N4m46Y7/uAcj
5u7ltfMgi40/pEyfgqgPcVqVAZ5S2FB4N74QbRlfHsfaX/fLX9S0Tna+Lm9hQ5KshzZVehkNLnS8
XL6quwS5N0yh6ObuqKxO7vXuhF6xFVDLNMranpF8FzYvocDwSs9HjxjYeY/VDZmKwjf10/xxnZRv
Q0NMiI/pqoUC+Vg+XW2TC3vuB+Gi2eor6+MV9Y0cqmCjvaafyK3FFD10i7/mpffhru23bWToZTBQ
Ak4CbeQNeNVp0J0dcdI+Tgds4LI93JLSW8BwdQ+0eDO04lu60VTvdnWXOpL+Fbf3ITNk4nTAWIrO
Mo55CeaEkO2KM9UI0J5KBo8CqDYYsn/MDSvvm25VJm4Ht/WAzAcOLFmmR2GpYVVyaEl1j0SoUjNy
TtaAPxxQfCDCs3HotUzutWX/pZ76qYlOVfdgbFMjdJq8NT4LmhBN1+DhJkRddvv97W733WHb6luj
2dLo3Ztk1nPhxz7M8em16+oh0hFNAlKFdgp0sNA7PiSdcS8wGxKQ7WQufmcPuXD1ibCIcqRdGpfF
AGcJT6AiWWRe7PY7COF1zg8bj1nNcFLssdNp2pMSEaLv5o47mCykeOSrI0bgUqFyYFYluI4cmTC3
nfsfVVWN7v/Kp/k0hVEiDOfBS7QW1FQ+2fbN2CYKZlblWuDDcqicZC7aqu7Kk+5VQYdJaE48gAck
ztKlUu6oWQZvPa679mKPBFUL8H2rrzNdIKEY1YQPk5B7fDejQmhxah32kwQMmOxxUgV9jxNKVU/g
fxErWM8mi+x/PKZEcLmZxdit8gx+llV/f2/t3+TKxBRPKi6ad3+o/StoGvhurZVyd7naPPi7AbnM
IWwzWDuLD3Ga8TMmiytjR4URkeWsWW1snmCm2XubgMDsiam0FgUEi8kJ0n2haR0DyqMG/hz6rZHW
Dug53bDfsZSWK5rmeBhCS5lGQF+qbpoI2MM5Xn2n5qSELcR69N9ne0NTSp5Uuf72zd3A5UClVR0P
KrWeGWg1C+UnvqlDoNOVAWpzuZZ7oK/9NrRKEWCZDIzVChPTTPMr8P6JNosGvODVgqKHTkE/tJJU
HLvv28Eox3yKuz3rwHhuBfmWd6ftOeut9LtHzRD0JYgkKBuIEbj1KlY1x8mxo1EHdxGSfblJ5NnX
upXmK1kc1J8q0T0c1lNTUyIPr8kQ5AyqiZN4jNyG+nSlxeHOjcabxULxGHrrf/74oDBC1HHAbFKr
MP+5Sxm4jNVCtuoxnhgnGG4hFANaNMxBrT5MIHFdXWiwO0YnQWBIPs+9K+XBw80O7nuyWexw8ePh
zZa/tOwuFR66mKR3VLANtICcPv1e8Sv3KH1xdy8c9gHva5IqFMSxufBFucMmOhH/++iaYHbUVyO8
xidel1PzcNC1SIVd7xzAX84IeAdaNkKwlNnWBpxYkOar4GIif4lolUkO+C0AkLOSEZsBxIqGTOzo
8Dr1eAkwrcfsF3e6U2uOEMxlFJrEg/UjCrnPv/VBjpsqSWRcFpGAs7kCGV8Y6X3m6PY6Yi1xWvtp
BNPj+wi1naxbTO12CRkiNZY3bcfjSa3C+RWG5504NDRR9xrWnL3SyDfQ2CytepSeoa5pARDsSg2d
kCRFRBsr3P9qM8iH9VhWy+0T075YQM3T1TWu7XZey18rq/4IJB1hDRrlOAY7TYFYJu9danGZWngD
nr3QHLhtuYmfl3bFno9CxlOqSCEN81FdZhp3Y/eQi0zFvUxokTGzR26IosZ6bus5wpBkcaCCcsjJ
cX1IWfL2mK1lq3QiSuoyj+ZapCSMinJ7aQ2fbtK8KdU50JzCyAEyK/3Zvgi637wa2bBpD7aP3g1o
NVC42Pkio4uLrngD5n1G5FRr+7SZsP/wqLVpjPSVMjylQLDshibAQ/KVXd3y9x8UoaeCC2oKqxMa
UnH99rlltv1QyrVPPy9ePAztO0OJCY/Wh1pjAbb5kKlcN2hAaoHX80OUwQy5+N+3oF8XORxKoUIh
Q8reHI5o/o/xhlZEFtiNMbqJSkyB2/MVwqcZ/pVEXNR7LCUxZaHrsvCTUrXcqJL2V6tXobasdib0
3eL/AmdzoiBEFnWzrZaFzfaC6v3BDtIwq5ihp+VRR3pnA0O/ocXraPJCTym12ynnlXEAd/F7IQYU
a1K9SK4X0ztUtRgSqs42lhUQ9KWW6At23H+bVhu/n2TlAXHTC+uAy2SLGitmWYF/nC5zbh8kKqB1
IM8SfIaFNZg5Tccs7HLCayWK37Ui3Ikf25cu7sC4vkOTxr76al3WB8NGmdOTEEqa611cXYcUShmH
qG2IcssPZW1Z6y7CXCLL7VTZIVNIIJACKN41NK/f15Ne1iN2mWF0BKsJpcXEvze+Mnvxo9D1TFaA
a+uX3DU4etD4swzv9CWEFrHada02zc+JI524ghJkpCHgoQwtt8LxrGqqt7SzOpwz26yWGU5sin9I
mYvZXK91vKnEOV8OpOOPPMrA/56p5u3+Y8okkRgm2aFmMeb/GWDRhWxY4vgE9t2oseVPqdGY1xW7
KUHnYVa3gx8t1oN1ji2nVyj3xSIIY4yMCED2ebnsgmZSk2Rj1/F03DCqV2t/uSL5X/J69UzPCNtk
LPKKX6IQO/8hilz1W5gKonZvrvjyXWN+y3jXne8uyKYhdaKDMRVOzCzDMLDzhLXywAIotvSljQlr
Hgq6GvAdHsGAA1z0L1QTCLdxerOsbU8Wq8qJ0aIZol5cF3vOKXsq7pHrgX9TdnmdM5X5tcJ85jkL
T5ri53Butjln+VxEoBs24jD5zvNDfvbjAt5A+ApiUCBYZe0evOS6Kl9Cf9GombQSMymOOOj1fjiX
rM7yc3oUvYjSEWo93rjPa6vwueQI+3fKRyfmRKDCkzINwPyzqY8Z6g5tkGqQCUvZQ6mGcNc4GqF4
gLXDoV9x9u9zGobmxZ1bwWFkD9AyvKeVmDYzpg0mjKs6G/dq78C+cjeFiIHwCKWTR8amwZPq/OjI
S0C+I4YH7KsR+HuF29FZv2TkpzvW9tHOOBFchK6O+KOeodYQk47uu4xllvvJ8WjJZxlBbQClENaQ
zqHqtMdweNbM80lJp9ol+h1yvx6VCtwjmGHGkyZYYucUpcZVcThr99EXK6d1cXsrU25zrxtw/EC6
/qMNak7vuc9TztiWkEhKKYK+tR7KyImFB0hBnLwgVL+GNa0QCwuaANaJMzBaSzu14lFwCg2AVLVt
X68MtqSVULxTZ9eVn+EF9NLVdDrqbBNEyfpUOW+Lbvn6BJj27fJb3TUQE+WGodnWjxCmel1SoO0P
9i1drzEZgCZ7YhkDW0GCnO7teO/10Fwo1LW1keJQN8+uyzm8KrZIZXogywN+AtAyW1vAEckK/51X
L5VHtIT7wKpVlOS9QkkZZASlVEV1QbXW9dnPbEZZFmvdRFERsvaYgwBLiFHLRKMxQV9ioLnwOJJu
ffIQzkFgzuHHnimgDHqBWGMLSq1fEzsPbife+DLf67rqUPAs0ypcBkG2RFDW+VkI5W1rGXVoGhiM
4gcFF0BW50JulJ5ENqEjRooVe4yqg61X3V9utcqcZGwoEPAELHM4uT9g3KmWHJhkJaCgQzpiSa3Q
DgnEk/50iIScN9VtHkj+pAiQPNZabsR9CnAY9UV4Os6KIp9NtLbcR8Eo5D4zk1gkDe3A4yT3QMFw
x0++5bA4HK10xNKTWvjndQ0tmeezPNwXkIvE3g72PlwQIaPtd50tH6cHcs+7Ld2yrWnmqwam4b2C
uPgTNLGvKgmkW+Q1kAiF/+EVTJVZPK9vYXTzsUnQgN02Xk5+PF6EQkz/jr3E7ickxIszgpZyLycA
g31yrMtteOLfUgapwKqLYC7Py1sDbJHNSSkx1rpAEzPZICtwTQV7eLWEjQGGrNF/EWjcMB4mF1Rz
iEDMmgI/CJVjeWkJySZ+4m19PikHwQbmUkbbpo72+snE2+UcTGmwFDlf/twjD3o+ymby6aiFeik2
637x4FBV6DQaZpgcU+RXho2FzSlNYbG2GXr9ZVM8WkmTsEvEO4I8oeZFNuAZKfjkhLigs1h24GTA
wet0nW0iPOJZVnuhaRV9Sy83KfGZUeWJZNbZIs/qLH6PKMYeOcAQbdPH89sRO8l1YfGai2i47/MC
FurxDCd/4Qca/fUIaPx2Iqrzo4lbCG4dSJl+sukUcSdi6fcikeoLswFm3T7mUSYzNNZ69/Vf4hQv
3j1AzgvXT6Zj4uMaGfZ1MRll86C1yVPpMbB2zqscWj3xpp6EHncE7ik8tXvcuyfibUPd+tX0ivDY
aSALcimk1hbX1HdLJAhfrv0AypaXy3FgOmILeISgA7v6qRDO4rh/Q8n2r/i2JcYSvRegRPv1zP7x
6MfiwGP0dhHySx5evo7OEbx67gI2LGaXT2ZvTX21wO7UeYCxGxnki/QSi5iOadGfv9sgl7JVk1fJ
tKru5QFwDJdVKsOJ8ZcMmZiwFjo//LHEMLw3S1LSdduI8XneXylQ02DofV1QsPV3GbpqYP8D3v7N
Qp6zESqt8/1hEFkt8m8DMXMKFQKG2qSBkJ16IXQogXX5WuzFvazxbk6ptI9qccv15QTBNZ8jugW+
/CbFYB6s9bor0XYQXqpCUs/rI/rkvCrfAzuR6D3DnAXJR/iBiyL8G3UpFtxUQTfI/Pc1Au9HVzvj
+kaGoDmbA4355/fEv6nbYpZrWqL7BulgUjtf4kfVlhr05uu2FS00NXmfta5VHpo/Smd39WfWAQpR
9MTCvnsCYfXrmvOCAda8NJFieitGsWyIY1UeaV7uZ40nrHLN1mjiEGFaiPweaI2nJvxhq9C8B6+8
4FgI0+F5QyvUvUSiTcbZ1an5gjcpm1OGNGVi4iX9HIyOewGYzRx3MbfAEguOCrNrfaR0F6xlbAkI
TqLT3Ak16xCosJPj5/U5ggLIMZ5xbzQZ7Z/sifEUtBqfhNOfBp9EtERKdtebgAB3xmyLwwMhQBvO
FjU2coHIUphg+VE98fpOjFYw/jxYqh2O76ih5tWRgQbJEUR9tVfaQmoYg/LaXMexPsl2PqzCD5hJ
30uZR3qShLVA2aLS+DV5YjwRjESe+yyNIa0oplRa3whz+JdjKZlbN/4pZABZvUowZEs4KYWgTC5U
enrbqBcyspcYsWRioBibKJF5a/wNdFht3tyFMYffgi/Oouxy8RASZjmkjHMqm4c4ju3Z5Wh45TMI
mQb20ZMjfKxRR4fgCq+86uqKnfxpoxKmw6VCQXoNj2nC8ubhieHnVBBoDcJXSOyfkJxlBNAv9Upt
hyymj4DsapC2548FdOij1Ce15x4uiudaXcMsP9f5GUFsCzfS8bR8AzrixI9Vvsy6xXNmA87UToot
FGbOYRjIRwtQEwhnfuEUcq7Irz8EJm2weXDUoTW5FvcxNGUxCk6IQ+svK3jCTjpywVp0DLWsJDtA
9oblZi14Odzh4N/aQM/OpXNj24YctLG7tZgDKgIDFuwVwIohmn7pMOJDAMeC5NfIXxFF8aCO4nnr
M7f0jT9e4DhI2v3XS3N/ANuDuFGKlh81K/xkbYHuGsKK9zLjKpytuCj1JICusrWfi+mwH+UxfQlA
Eq24t3zDd9YSoCvzWanNT81Gz8x+0Pgt6DHfgyxbTTaGBJoRvcRPdCSGzL6yuc1/P61lrD0+cQn3
gZXnGyo7NU25m7Aqte6rlBao5xaXhWdGkoZcSN6A4KP5hWyQzeEJlR5W8OnwZ8WnnFFb8IrorTU5
1rD6aXzoM3AmXOjegLGHvkdBFnmmhAG+q60ard+wPncbrKU8M1zFSV3UdNTHBWHakH0KbuBuRDxj
Lwy97DMI0L43eM2mxYDnVrtp9kREVcjFOsfkNXAcZXEhCqGiuXO3ubDEDHj7u+WmfYE3qKL+NziT
LNqRnGdH2zpECruxnr0fjft0WOGLHfA6FuwyHg9gEthngkhR5DkCr1ZctkHcx7PN7x4OWgac+8Ks
x5XNtLstp9svLX4VlNo5WZW5vPDWbLIGTHrYSSUutC5oG5O9ZKJKC3mi3j1fOC+67rgZ/nIAq1tQ
vmLAunqMICvrIs400MzDJudqr0NYuHWQO5ZsK9waBEz7VE00jS2fMhfZdC8HjYTlzKCjxTfLOkTn
WsLLn3yS594nztcbyGeWHfVVLbDkW7Ab2/vykoBfCSbnLerC2g/CaXSyzo3r8ttSTRmv9QnbEGy0
W2Cdn1FS/FHBTATr081F4ZZyuzxWabEMyOQ6hj8OXP34YtMHEKxjeS0ZL4M8TI576cP3eN9xkmWD
5EAs3siUg2j3V0SEgxbD/0sE7p7ZwVN/4NvAEeuPgHGTXpmseopd+WYdh4ghV6TYdOVioXPo/2br
nnWcqqIJEkdTNewK8Q4ITkRGC8qLbASmT4SeWMKnmivx8gz0BJExtSijOBMAk36JyH/98mFJian3
TR58ijIs7NEb0xHuku7r0OSLbzJs+YzwUSIIC1cMvixh8epTrhw9GRsB4FkDOsA/8NdPQRNWKhVk
ILsdRY9OhiWeRGSPN0ke3PYa64fYZd4EOlLVLCkMFHoOXuEsxenTDj6jl8Zj3E/qDeYkdkQj/Orh
th/1tEP7zTWs1hHK76FOj3+eQ0ukTc8uAZuTfSHv2YaGpkeN53QQoX4SlvxESFjS8s29ixFuBhAT
EDcpcmvmIed7f0vfq6vPZsvKImYOnqixDVN/CVPRhMFeGpxL2k7TjmvHmoP10WnftwdCHL3FA1qN
ATcqDWeVYqqfNd29I5vPmF+5LKNOGXcUQrNX05KCrV5rSXMChFSE2g0johWC1ydHGgyaD9Hj3ilO
6HqlT777ojd2amHBpk13IUFBrVtxUIrBvyT3ipPGDYr6PZg26T4uGOGQrdKCCNo8BCGoJhzxfIy0
3AALa+pU01tLc5/VjTKlmYLXQFYqepDU61pCQbyYO2HeQHV23JmAbp31NMEwRQai0PyF8w3qv8ED
5aU7I+e7xR5miNdm3foAdMFU5jfM7B7nHnIeMvenLi6pUBuzhAE8vDePp+9ZF4WukWKNoQ7/tlny
uO+rms7phY7IfWKJ7aOPZJnHhUHZwRNGwE/+Ucoh6DuPu+Jest+NDjIUz0+Yd8NSybeI/s4eahG3
vb48KqqHfxacBNaQppCVXQFpoERMhJx5d2wif1oUdZLW3ibQIa5/AXHLLc2oqdW6w+fdE7Fy587u
V2GzZVc2pe3ncB4RFysG7iAwA5BtVWLe61DRJ61yEjSo/vY5TseGqP2wAUgIyXgEjm9xLaPSnFcu
ENCi/UZVHGkldaH0kINNBeuM4ebU1JASFiQZiqOB0JXYuQhDyuN3aT+U290TsqgCINe/8R8eMOrv
KY9/I1teKOdhWMvDYxK3xCMTyjA1YlzdAcIaEqHMSuV8/9T9zffwbKTgH0KWCvYdG0H8i5P/sC8U
tgkA98yfNQ9Y7LGqtmnq8aIs/mz7NxMMPlUo4KPQ2GFPMQGLn0mwdiTwkFDAhWgOfrmbjCEGQqya
vuND7ufU0O5O403Trt+dIOvg2UHbCnmT65OjZCvuhXd/ihbDpJEQMFgz3qm8wWd2AfefN5WeB9Qv
zK25tohvN45bLzyhp/nhvlqWfYWAPmE/NoNmN4u7aUqE+KV/zvr5BXE2ZKMXaidcf7HOyV9wlLb0
wttx+Y5eDurjGCTlpN+MJYGpuZsF+K8AFJTwJfy1WgKBe+vjfGSRE8Tt1p7ZWgwEZmfaG7urFFjw
e0pCvqvMXE8/zmr+XMgXYZycK/lknYiITaw3MKEJzNbvcqHNB6aIQW4y50WVkPZ5TBa7k7esmzQn
5xjHLif1PNS6OnFxD+hFpEBEzUKKBjbHUTIH9+b6snwKoTGbAJ3ObP3vpMRUYWtkB9KyuHEe8Fuo
WpwOcTmCXGDS4nGd7syCqCTdrVN0cWixUrax3/39PztRHHqrsEecx4c4hZ3j86Gel3fMOYewCF/R
vTQhQ1W/F6XgkyyipV865pyEf5fbED1r3E0MahNNsr1g1D1jXOjvtuLFaoJsoDPFpQhr2eimSr42
fGFhynpoaYgakefupD/Giwd9r9n8F9qXrXqp2zZBVKJWjYi+PdiSHuLTJ6TgYJYCdMx1Tz4hopqx
Psp5d8APAC6HtIbcgrh2TBiw7QK2/i8I1611T4r3BT7+XN7CR5XrUwuQe6TWutfJuY7NYWve97e0
iCyiyKHFGbjM4ZflvC9ChNiZbg+ILm3EIvbKf2sRM2xlYWZW3L1poXzGiWmODT2eAndGN9sYDzvt
xrf5JVDyaqCNns9KUkjtxxDGdSpbmK7CZO2/e3zsNfgOMh2xqfJ/1pJno5Lemdn2NugCaQou/VBh
2M6gwdVl/QeJzUsFfh+rvDZEa4gGbE9PdS62rJrJQnPFg7CEt83MN8PDY420hVjWlUUERSYF3hJk
7fSbYlIxQagvT2l24OaZ2vDsiR28rw7eMGWlsqtohUqf6I7ZnmzSYj7T/CTCzvdesIxUpmaCEE/+
MrJtUg6pwhvbSrzgj5Qp6NWcXzLC0sOeO8Q6tgcLP2eqUMOuPsYtn4KaUNHcjpPBVrh6AFtrneTx
v3obPriHOXry+LbrBb1G2rn5UiUzXc9yX7qdd1I7gk6EYsf7nEp6GjpOBA1LoVnB27Ga8TNF8FVM
7sna3IpyoBY2uBr5j5Qs1+EdDa7tBuJFCDI4aBwZayApWaOfAwNNJb3/FwDJQJYCnPWpl3Mc2p9x
ezicWNbmZN5//qLBiAJvYnVJbETMGWrVU9mJ49gtjjVDKEB6H28IKl1Ajef3S49nAE9Agdol0enP
ZF1nQEaND79MpBw/c9VuKLSZ8OQPXzX/Ypkpa594meE/RoiVDY28iFlORSpX6nauPKaZfslMuK2L
q8xkQh3bpwxHuzbkzYp5QanfMl+7g2+L454g+keSuiAPgIoqUdsbEIHeb9zf2cu4D9p2BR1SOkzO
M6VYISKnPf2DQj9nmBRMXaYfQAub7lg1m1yU3LApuJP9QGz7sSFCoWcvmOpBiEk6wOr1L8od0hMe
UmWFzc5ITzhkHtG3RkfpNghPDgJMiluY8bLbTNrgF9BiQJqsuCPUKAYSFqOOApNFAYItsxX/hntV
95V+Pf7tFfiRZLZCLJyo7U4tAX/hihECcriTR8RU0n0w1vyx0W/EkajgshDWH43YQtioFOOrx2Re
J8M6hrUubPLq8REO9jn0ZBPjn4ar5+4H0JchBrU6BkqEo1h8Wf2ti5hIC8LdZEeXnclvX9ErKn8e
Qgs8RiDp8ah7bqiWNAkoaRmew9bLycDtWAOkp3Sd9HqdMgSLSJaxedpFtcTYSDK0WSUOAal2Prqw
RPU6UnlFNGoZ1GLPs3xP88uuv/8AyCKocOjT2qA1IGylzHd/WgkMjB3Qq1gMP6H/h5geQ9lzIfIo
CA/JycHsVaCnbscYpw3bUuDoxFwRN5TfQ8mlrw5u3uQ3G1Cc8x3ZIM7dhDHVYcqf5x1cDW8uU+Yg
MpePlDL38K6DiLeYG678VPuwYLr5fzQolzxnJ9Z9V6Jz2p5/sgwTnzU+P2dzUMr9fKgpml5Ywx2H
0Yaw75aV5g07GeG2NeVU9hF5sDrlDNXsPv2LrVoNdzJWLQJc3Fn+BCbRSdAH06cois/XovBWb6Y3
d/TmLndvUHexhMpaVGbA4GpRiEExPGLAmZTaTNKXmPLeZFng0WGO1uY4ZqlQB0f9kgD4RupT2x8i
tW3fiT1eAomhgD/ayyyC/zJmhrBIBrM7gaof4BhNzWyJr4K+YB2z/glwcGwFlr2IxGDjpfXJER2H
gxD4ACodNv64IoIZm6rKAQGyUy4FDVjWeEx5QE9V6l7mLquQKLpG0w6Eq1OL8aFelfz2y9kao2oZ
eH7SVZN0DMCOVGQCNzW8gKzBlnZlkKAx9utfgfgsT70xh75CQvUPaBVrMZaRqd35wB95UduGqc91
mbNQj0Zafnj+zSvMh0rn02+l9XPhcegUTlM8swYFmkuCEAWyKwbiVhWekgKaC3AWYLA4JAeBgWRX
1f0z8pL3I4d2duoY05MNJONrzN19iPai9IUBUdcDfTYxCupPWqjemCtne8KCrnxC/+NJ4UmPuTpt
8+19SSSuh6c1wI9UC0IYL5wKEuVHC71eh3LcdC7GkqYhVHVPRmMFcfg45GEhRMDzqyywPjUYmq5g
7QH9Nl5b9nuAilbJnSYiS10OTosQUL3bzZMOt9447ekcq5nmKIQfUvCAL5aQ7Uqs8nKIupV1U1Fo
L7iZYbSpmu5nkJUwfSbxeoyTQrzGQ3q1vgqNYkQAE7bUN2vGyEVVqjUoP0IObndKRn+XtsWr2YOf
2ws/h8RQJ5mOPHraHApJPRvBeJ0ab57Gb9iPqlIMPWD5mri0tWwnVJKh+LQ/Qhg2h5XGTerBk0Jp
6Kv4tyP04ctDBMsyW83Yndp8nuqzFFqBOYnmicy+X8sxPYb024r8er0TSoxUSNiaSVqhHsmTcf29
6VoGijKIMGNuZ9W1MfMFx5ThW+LW/KvLJOtSg59BGsvaEeEBTIxEr+tINdPUP5ccnMEwHsjJ21su
pLnYjwzebdRfjIuZ/gmQ3Ck6WRF3yPVDvVInHHseFWOXGlf5ATUTNrrjRaDTS9EzrTrVEKj7hrjm
xe+PVIB5jPgnKBl8xOycDWRZMy3gDYjp12Z5XgjNqt9uwoA57rPK/882dyew1ls7MXbEOSvXmzrV
kJ2wWX2He08tLqKsJhR9K1YELE5P8zfGtiEcdSbJpBTOLdtV/gbNl8hiCDPLdkdxuURStnUYtKbn
xnR2PLjvhxNPoRW/yz3a7X9PGVKFGXQB8G4gs6hbF7qQzhQHF/8SMGAVFHEKm91Nbn9K0xTJm4pz
owDXwScJTtl3g6oR3dB0c4NFtTP2UheEQ5CJbVIQeHk8qC3XU9xN0mU2T6ZOim+9ZVapSsAfAxjB
lrmvebeUZPBCkH/D+uQbDome+skYMR0OYHyTdnjyvPqYZ5OiEUEefecEIRdOFA2hZwM+VF/51i97
IewrxAtKTOm8ZIakBjJCTEUtJAu1Svb9WzHpXFMbRdfrtG0fxHq78PBh60Urb0kqvaiHJbZX0trC
rBM9zIcyTsjIRLI5QXwbaUVELCqPkvVb3RzCYwJwy85hyAOsxguTmHyuMCsA5ThYKWqTieHkL4a+
kPvzvVMa2Iz2EWo94qBLY/kzc6flSw9foyhIa+UZK64nnyxQAyOgupEpVuAIG0y1RnTaDqu/voXM
gFhDsIWBewBNNCrQI4fF9SaopVyA+BxKq8n/FvbRh0Ksj4+a6MFDbZTvO9ZzTtYLJYP2+h8KlPQB
QZudzvctVRrek/Knjh/2n2va/zkEqvhCwPCtQQDUWdSt3CUDlfaSuV+a6F3+QsYVbrf+gnXOlD3F
beq7JzzcUKTkyCKYHaSasinkjW+XkfRWdTZ9Izp/bXgwoemaNf5LLUXq2tRvGoqlSVOtFCF+UYI/
b9mpt8P8DEXpDZueCJmd/HgWTbrHB6sFOHCUulZ985byYkJaMErY/ye2QJtNo2fT0/Ryb+gG48oO
owhBBXyhsc9SxlcehMZFoGdFipzLBJTcv1X6j6BRTdRBvFqj16YhK0IyriueSW/Wp/Gmf8iwTuq/
i39htIAkYrVQkwwzDvy5MAA6nJT+sa/GOTxM86ZGgt8ieu08cDdjk1IKTXjIJgWPimmJZ/8f8GgE
VOqWRWOfUXxgEpnuC6N0CoNfiD4le7BgXjEbQuUeRYEl61YYmDXZ7pV2f84D5ZMPhvwl3XDGsvqw
NTcxq+BLlTAGlgFKSi2AW6iNEE32AelOhdNyTtAFkyrdDW/1YnFc7TG6N34LQb40WTS1RxmaoKVz
4JPHEIig/9S5/f4Z5MhfT9hcJZDJkQs1tYjeGw2Ps0HLvt+dKojxM9YNeBm6YK7+ydl7ue391O99
3DTcP5WBeo33tXv845Fh2CVQwOkwIpfQsWXJsJpXmk80KkMje7xbheWON2ujSTA/3OPC023gcgRY
E9BmgQOG+orqnWu9oa3X7TcX9AB/B16n6aj4PtxwC6roa2nzy7We36XnjLOIobOMmoDwpk2a/bzn
SqvTEqmduknVixS3oeeNdaOleMzkEOCGtV0rSI+UBtlyEN64ymT5Wq1NfyCzIzwEXx9unWGi3Oa7
8y5QCDMioiYMJJNPqZxBQERYR/kdJZCVWEXiqAPpdLXPd4GbLoXb7u/p1HYTCghtUjcBwqYUmuSR
ppCFU0IkFCBOlNTMa4YnoCqnjzBEPqu0uaGa9wZCUQucjxv5IzQlvk8SCQumVNvvtSKMOyRMLp+Z
7pJq/UjWzLLcqbw1PktSjQ5p97oLg69VHt2ALdG+Ff1VzDIAuTbI5qWEB/nonSBGWS37RQ/nqZAZ
XHWGi45+dAHDK1OZj7NGfTSfR7+Y+SsiXTVIYdgBo2sY7sHBiUqIBiPVuzytEPFvKKGN2NjXfEu1
tft7joFQ1nYG+F7psGYQQxlDJ2RyEIUyQQdCa542YKp9LXjGoewYwpHefjRCkTGn3SY8o3dtAKlY
E4J5LRYV+voUyI4iX/YCznIt8EsST+fpT/0NtkpCUjSzYWCPadXClT0mDB4/PbLUnrpy7X5R3srs
vxpG32F3tFlTY2gik48x12zDgz1IVumb/s/9HTCt/P2IXx8mZ4h+5DlBIlNvnq65Aiu/qj2pfM3h
GTz5sJZDrTRPoUK9oU/0Mfw7UKxSMjLEBL7ZfEngssZZtu6pS4dHRWWgctioDgc7a9VmPeVp8QkP
efoFV+m60P5VOE072HarPiu5rx3cxM9Jo3WVC5PfOUbow1xEFT/XzK/yWBWuNKzPU53P0eq0t1C/
X6Xzcu+1vQUVxSqIEUP99jVn4zntUA41W57ji7f4St6rxmigzaJDSooSnPt3IQlWRgKbxhYIMurw
W87pHgoKnKmkPEAJ4PniqBFFEISx4VcobYdJdl6fnnl+RJZ/41Tp0xmCuBYbv7R2SKSlfPd0jFRJ
TXlpIYAJ2bwUyLb4oWrZjlWreZewP53B28eJS/atxeAQLZ423UmcL58EyQ2zaTYD9mT0OPac886A
550O1MWGIOMA+DEImqzP0Q3ehQNhOFzym5EompgspxbdvOAbEg/foirnrWQMWFlDnm9f7Knb/POy
mZeByZBj29IosafhRBaXDY9A1yC/5AvoPUXBeJRhJzBCuDk46x2sEfmn+kaxmYdUVZYXf7GmUaCe
2fNayfMPwyzeiYFDOmwmD0jVzsJy8ly7vZaz6L9FtJBoSz/hpvcN8NB6/U6Woa/mSjSnFnuft5ap
Eiqigw0kxvmx7uSOFnQpdWpvPhtnEQrF87CaNX9P8NwD+zq9Gy4QgwVCfELsIl1v1qU3SaqoiPdO
RW3a1mU68xEizU5qFMiLdCElC7Az7Yoiv2m9uo0ayh9G76qgfGiwjg171moAVoxHM9p9nzWSHJUa
u9sVlbmgrECDxOhm3r51SEgtsiaRwTSpXy56s/fcC3kPo5Dtn6UNBogZu7fKKTL2hWU+Vyw44f2S
0MimAXndpHrlLpP11x+6efnvuenoBXPSScluseUbqzRILeC2iQk44pxgEa1cc0DFqtUFRV6O8dNx
WOWJqoQcsJ8t+mDWWc1CmEEIvvMD4OIjPWvEkAknpmwYd36o59REJqkdYSr/fYlBDJVnfRPRAiQg
tGe8a2Tcy785MGjv7HEQCwVQKEUKo0IVEAmU4FAIEAdj1wiahwNwLF/3AyNm5DFt3Jcpe9z8DhVO
5WXIw2EbG81ttqhTJQofzPofojp+avzbkFEzCbXukmgeELyh7R+Bvz5L3eqRc63PsajeJL9HFAYM
+QPoywZPDqapeH38n12+W6S0b4T8D9PHytv1JHvc6An/MMjkkAYx5fLPiZkFGw2xniLhAi9Iq6N0
SrK0VOElC/C+gWQb5OVTrXsS2aCjkzSbwbKMGYc11RyAxjnCnGSluCx8F208p9ZKSBWKvpxCSS+1
p9C8J3x7p8gQr8LGdtZW1iqU7ZmcX3sE7WGyKK8DG4Kf/4Ixtwc7P/YoMxwHQ6L+qwML4Hsdyh0/
raFDEhy4AI5YUWQEJg3hfYRbt/0Un7Zn5XdH5h8T6XcmHB7s/RAp8lMtrlhhjvAjoH1xWVg05Xq9
KBtJUCgheKd0AU262vkkbxheAU40BhHB4uWOcTAD73C5GaTSxDkYcIyQ3LjsGjU+aro+a5Vgumpa
0vq3AY4mknTFDY8piA76q540h/9o8x+9NUnfEPdmeF9+re5TpfqbI4GCId5MlYdYZEb603SKex0i
4Y8a6TJ9hykwkmBBMnF2Cp9adEcIHbn20UHXls1BeMzFsKJq43tWINBrDlUdiu6AKWBXYOpIM2hW
N1tPTvKTIuwy3uKuauJsU6wo+FFAgQBHvPlvMfS5Tu/2K+NdnOVzYCE+44W9B4Q6iADoTmVRxHKZ
aZBf6/IMkmxeWb6NsJLNut6TpDUvpoZbNPYLBVmQPNH4TGmkePKQly2R6/bDrBoXkvdihMaxz0zD
twxE4zXWGs0++EBP0reKSNSMO44jV0duqoVKlPlt0eoceC337M2WZJe58Z9HqSq8m2O+zG89Asji
q9aOtum51yGV1e6zXAjmctkSVDSm03ebHS90UpSowbKBdVLP4i1jeLyLgJsvp3cU0uuJCXj3cMAH
H1wKCbQD9YwVJx+IoZkPiGU1PLRKOrmvMrewh8iqPts+64/evj6mheCoF/ZDHYzS91q881wyoJzh
SvqMecnBinjxKtrWs39XCTIWYemfexDkkdk/EruO+fx8vpH3rgLU5M1x73gGAzFEByAqGoP9+z1r
jPTUD1fn+POQ772/BepmOE5nHGZoIvpT6dr0pM3qUbo9sabm//+7lB9Qos+gowP8MC937IGgW8y1
Qx9Jeujy/am52QEzkvhBb643nJi+s6EENo567Bsd2taHkygiZxq+S8SZa4Bj49zDKMJeUaZhYkQd
f5ALR2yW8jy7uljDW/mIr+2Ikvh219DmW4kcn3qE90wP73L8MJ4PmN26ZDQ6f6lZbC116i1OM86T
QuDZKgjKNEjt0yXOx52QfwiKQqJx25H9fxHEyM0SGcdjUuhE5mXRUyPcJrcbTLxhd2jqSHmOTAhY
oVvY6FHTH8sThJ8a/PRO9oJz0nP6ZW8W6jio7s3avbJ1xU/VbMnvE3VtcgIbWFSJrLW/c9l5L7pu
bnY+HHx4IA4+PD/+HtXgwYGLOLPaZZTLqHzQ2AY1E/QDwZk5CY/Js2sRsNHrYzsdq1W3ge/d6dFw
gSwOF/p3FeN2Iw4CDTa9/+JIB4Vwe6NEPYiDNVdhkUiGOJrI1A9i0/ZzL1as70uQQ3VQofj5BzxL
kZVPefiONwBnIFNqdNFvR/64RM3E6GJfyE52/8uwS6/oVC/RAGPIcb7B3K3aNUuthgwwDBI6ixqm
SXb6B6g4hx2MlPr45COulYgVRpAEbopsBVU4O/O4k23i1V703sEn53Olh3CVBbGmNC3yiykkm6Xc
GVKjxW6Vf/h33iHIr9IpDLe3+4mKZdGI45zww876blYJF0rp1NSCfbdb51yQVL8cBfxezHHLYZGz
3mEZCdEW8u2nLXZ5f/EnQ9l09oBHWH0QxkIp3XDAL8mIou1lVh/oE3futlzGciIADeKXoBCMvbQ5
EbOSRDgelkS4Xy1Ofz9pKiD/bFuYHazpRoz7ChPZAKUEBEAhnjzwEvg13ujHV8ZADwZ9c5k0SaYB
24QdQa6A+nN0sFZYgoJNomPeHQAZ8aNGVh4p6hw+oBPwQIBFVoM9yblP0l7k+YhtO7kDmNnmHW3U
szFnD+ufRGLa3BfctMYuBfSRUe9tfXM70P3r0VnJ5SiUuN78vUzMInnQd/P9v6UEHg2590BXtddT
wcwxleAsnvHck5wKFSYT1AT/GhHFkupU+dpOLFXus/6bbw15BJgsW9QBNvRnn1YFg32xesxmVwK2
5CRqg0Rkp6MEEW0fCfOoe4t4cecJgPbgVPrYyS4flH9hf8BpNd8hhxwGLfnW6VAELwt1QYbcgwQj
Crd+jd7o29LhXOrIln4A1Ab6YLK9KXK6SOG/1DrdG2asfrsg4ZngBSKBSol3ZAzi//es4y84Rgjx
km0tqbRSsxnW9o8IBPjq2pOqx7WGwtjCzrSGkjBS36aC+pQ4AgCUAu9oNFqt10R0a5H8hVGIj6nK
vjcA4REUk5zCdO1P5dXaH8cXa+wg6d7zRH/2Qh70OHrLJ5VZwknrZ1c3yjHv1rXhSAkTJlGiosEJ
c1vEJDePNlw5880/qkBhnlSKzjP40NWtBPM2aSCNw/IyvCGcPHx/nnFqC8qGs3FdWkUFCWYQ5yzm
GsFj/8cVc8gqcUbSH4/ZNtJXIpBjXU8F38GlUBiL0Js5yNl2YjuJsRfCkYj52/nZT+fPNHJwTdBc
aFH7LFBA4AkkUFMDAZEAE1ry0/BC2k2h9APxj6SB1bJLmwuW9LtR83fjHN4rVdQb41q5US7MI0+R
XIOp6A+iJsfQdNgcxISxOxpHoIBSjW9YoRuHErv7PfVXOVZBDSF9W/uP8OOAHlNY24krtrXQA6rm
pA0bKxpjVSL+mrlB+9qOBdiAxqS1cukITsT0t0hC2aOe60rMNKsNAmCYJsSM9sFrhBMTTqAYvqBN
W/xrFrYLz7dqmRpWnY2g8OaocLzNiKL1zPJU/OhSHzjQD8e1EYQfFrHIuZ1gSbRBMLWOi2seZ80P
Rt2fpVGythufio3rSb4ko6rwalnjT02x9+fQA2a8plS8wAsqB7hcTLFW8nNiPr0UsWJoJknmnDxJ
mlu8tiEOPIhUedOC5rrrp3AHn/8UfGudbIb6g9oO2GGsaXPupVS2wpB805+4hbYoOx0KVBLrRwcK
xkc8PmlagQtlxaQbdTeE7/rkFzfeFODFa5z89hBopdEfwrydck6zZ0jnCuNnU6EjYPIFIQP02dZM
2e6De1QYAEFFX/s5Eo+AYqNJgc3T9V4I8KY6lV2jb9lQJDXkFKq6NEXHaADHvW6LCONdFwrWufXQ
AIYSmDMtsCDSTlwV9VSJsRsob0YH0otyoaooxpD2gzkG9sDv1Av8yY5TvkrX48h5jbex2TKpiqEz
WGdke+y8uwt/3bBpinGUke1RLvQi/cO+mYYTPy7s8A7YdG0NCrgnsQa8Rip0voV/+l7XY1zA10KJ
bJBkelLDUyvSCE2cn5kVBIjQcrHj0yapVfaZyCsh27ZokRDIgAm/Fz9weNfYe4FAwozLVZhl4HEK
wnQ/337lNXFrZ7LO8e31CbQ9Hqt1h7YcaIc6Sxi8MvuqVcYcaKf4R3u1myP3N7pX5tDAGS0FnNyq
BcQGTW0gqHUlZ1WKLy0fY/OHSLP/W9rErigWMk64QDDdNXhD1PYpQP0O1SnYT7ubo1jfERBxMBO4
xVXYLnSboUK8VzJkr+Kvw9RHu99BkEPUNJpfbIlw9OUm26PC3yXSUyqckVVszR+FtxG+M2HPTHEb
40F8fkFAqbnoFZN0FELo/b+ntNh+SUYuCA8U4iDMUfI54OAUz/boMbBn9gvv4W6MgZEhPmcrXD1L
lMcmaNE+tZvD29ApISZIsuSHkr9WWOwLFjEmRe3cFHd6sg3fG0CjdA3Gkv+/pBady8jn8/q94SFZ
by442PlSPA4V1OixJR08zBrTb5RlKqLEZtY0KTaE6j3YKaRKTypxKckz94DZf7nsAdGGqLqYBh49
5lkg1F1KA0vkoE91tHT7tFrm+ULNIEDLOO4pgqQwcyY972mAcNXxoZ1H7yKqjBC1y5Uud915NAPm
T/K02PT2EoogPdt8XbvHPjkj9m5b9j2zKPL65wXyMFDcvoB5iRPj7fd2w2rEwKupINxzB203wiAN
g1TisLmFPm0PYcIJjTQuYQHhpiAclDf5v4lm7YobvSVRfP9AjSFNG0lxkCtCLmModw7MbGPSI+6N
6j8kqNWl5UBgwFd9l9ySs8y4CBV9D2i1HFbidIPVXKQS4FPJvgfLsiJTozs6pbfT2xd3UyOjtbq8
hUtzEb5zH0vMeYhQx/c7hHzgUO0scTd+6SNjmYG6LLZd0E9UtKOrv7oTe9usnwM756XFRtnK4F47
YSyZlXtNZz747gNUIVtD6nxA6fCdkqNGlLO8me2vR/gUdHMBEalIcCt7jTXngmbPAMGn36rQSmUC
RLV0MtKKpejbnD2bQlFZ2RGUjVPKhbklV4BZeUENrl9nErfvmY37pJnT9dOLQ9u2F6OvZAHP/IxM
o9fhn3Yk7YBB2C41EQQ4mi94G6LygD+Y9RAsY6ygaOPa+XRbgNdTccr6yr0KtnW59J21SG1q9nuV
Fn5ed/F1MSgaMgYP43aR1EFmLeDiQi6KKhcyG2K85lb5+5c5e/dsDMZ9YsHGdIy7ffPkK7jSNEMh
dDafyIlxCjzNcsjlriIuHQylLs5imAHJHvT1vl9qezb7j7KY761XpzvWwJhTMy8E6D01noLtgl6x
B/8PtjYwKG5aIXoiRKOBarYuWZlfhLCfopa36CiJNG5d1Kl8Yhc0HnYCyp0VkCyWKWFGH/nA4H0p
dqeiIL6PccI6vcZYDT0Ggr/RSKDHn7vBX3cuYA2KHSyOvtbdTCdoDGjCBxU2IWCQAGtIWvh8JzAW
3SX2/1fAzqvpaEnnEfBETAit2xHUzPVVyzNtyotcOtSFyBSz//wXIcf5SLq2lk4d9E1TmtihI8Cx
UcxTSCsVTjTthCOyKV8/yffYb/07GO3Nfqd3wMt0EYpCh/TGUq/OmanJfv7Z++9a1+tFWhP/wJr2
36IC6URDAi/1tYQdjZAEPW97OINBF56rS3Sy2ZHlHZ4Ooc/NZCf4bs0fFL+t+5NtwC3UhZ/vfQm2
Ni85qfz6ecRVTv7yJwVdKRRiDkq+MD0/2S9A4kmbT0cDxIoY1ytLU17a0dBc3F56bHJvkaviae1a
hts0Z8n3INQCmxHAr5AcSxbMzHCxr6kNEPTYsd/n8rHgT+RzTL4IP7bTiOVuLNA/AWqf6asZ/Im3
i8Sqfjwwlr9CKBOs0gCJnJXuHxoULl7nKgMfQ98JrtN7C2zqrgQlgxhI5/8S2bxLrHF7XIfoSevD
asre0Mdmz5ZoUycj0v+ArEf0EtjbhLRGNuMOADHY9GYQnZgHqRxaEHNSu2l0ux1MgUsgBjq01JTP
w2QvpgcSGLf6iehGt1y2NqMRYE6RH0j2MdeIj4+yQcCsVSMxCL1wygJ5Bn+0/D0hevg1eHySP+Wi
vD1GWN8YK/w7YOX7zRrugp140qM07+QNr5+Iox6SenblSmVNKHJf8mrvNZ/N187SZ9ZHSGayOC9p
mPStsYTNiePt940xDiAh8MHzwebGE+g7X1UFqEJ68Rdicb/ETB3v/PNilFielZ9isIBm+euIZzaQ
NU4wJXwq+87Z9X1uwRhFWSVO+meGT9ESLxXSlqFlGJXGgp4mI+KKnxFFcOj9ijn3CXJ3MnZbrhWd
DAiXlrW8vUCRhyFCLdlzpGUYecqqljGybHgCP93pHu2Xcuc0giECcat3fRfJJKWSSiTG6gIkz4c2
e9Wn8KZit4SjFh25zGQ9lO0OR9yc5qpexYcwcYpMUK2fHGWgtX569Tip709z4kwtm3nYGXg+tgpa
Mm+ojbMG1kl34z2VaVXpZi4b/Smsb8VykJ5ewpGntL86oeETTRAxxZlsMd6vseiKBC/tif3oWCu9
9NgOfSADr+u772PeOJeR5HdvxWHArrj78QFhcU101bVrgoMRVhj+33PyPafD0pGpgsXvfWxw+qWo
tpuf0X539FHjSF5D/iTqKuasrtA/Nm58fyxoZZ9USkkTVMWD+U0IbFZ6DCS7LOa8rjf8PXP4+JwN
chrPONdVtXcel/fs8LjcbqxrU2V423/VdY0oSN/3a66+/qvKiMAisMFj1DF+7yCnRgkM3s9BhvNz
IJ+LYMbouIi3DbAQhYWwZUY2fCARMtflbyiAZdm6Kw8UVNlmGONDg4xcOpN2q5P9POFyVcpdyPPi
kpKIdvaxnqlXGdNcvQKBELgj0PxF76vcU6ORJDyJFGBCURsYGRWrONCxg2ys7zlJxK0B5eU/9ilv
QVhBWI8+CAIJYJctrBv05yeJwDVIp4Irff0KdgMpB6srGTd6hOnjg0FSAgApg0253Ao4qjEOpJbl
/HXu31Of3SusNe1VGZk0rlIfsaFSNNa8R+MVoENYaRkKYnBiP6xZpeBc/U/d4U6Rel7zqP2OdV/+
cLb4/TbM2pqQgoU2q9BX+ArnqNh3uNLetzE4K+6zhGc42ieGXodJat00kvcec1kOPABpvROfVICS
wLd8LKSAsLHJGQ0POMG5rYJu4CNcg3DjPWiz6lUy+XyQKX7vANvWJUFkEjNnsNJZkKAxP8FmhMnm
WGIt1Tm/FadF3vHffANw09GaVbtm5QzORzL+WdgphW4qZ1hUfd5+tf9Ui1CzNRxvwqkKTnDf9mV1
mJd1uEDWmnmgZj++LHPP32wAC5UqmoKksFDtaPn388DgOw3f80jpakOSh9BEcikbQhNszniz5oHt
SpmqLfh23uEulP2Uy3XbOodEaEuUAwQBUSp+1XyARaY1udUzSnnKWB9C8E+wFmHUf5H3wKZj+wFo
QoxGEZZMPAQsUx3pAHJWunQd2R1cPmF+h8Wf3NbrW0aQxhpn1RPqN0Q1AyqiRLLE9+d4NZGwrg9A
2pIBdZjQ5YZX5Up44AOHwo8C084sVMREtB2ITBO+llf/H4Ygk1ySU/8EHxtOAt9znPL6ODazeOGa
jB7M4yNl9/bGie0Lp8wOVI4It2VdK9mjoqMl8LJuBMWuLeWwO+GJg3yeBZCINTq4A1phiStibq1K
rQOwSt7QtDkKgRzV4Ekjn/07vG5ScwyWy9xeHRDCZ/y8fpur/9nigaATmTkTPhwh8GLOM2FDFqUZ
Fv/M4sihif4MvFfxDUPWZmthg9QD078SHT9z2ubcHwEgI7Hu6yw7sa9tXxAUwQRsA/ugXC67hL6D
c3v+xrTztl87EoyxsEv6YmWm5sMe8+KWSgpzrd5DfdZ6OjijyybnMlJ+uQ/9TM+PVWtPZer1aX1O
E1iibWV7YKStBNTwtn0aorz4Dx5RNVfMRcRfYIQn6ECRRuoJq3D52YoL0kPaAWToscsnDL73bmCs
KApSdldcsRlX/9Nw2y2TJIEQ/L4D8Uby24vy9OXMKki3pBgzfciCb7fLOLX7QNn9ZF+fmd6ULwiS
js6kkHwr9ZdP28iwOcP2aqy5tJeSEZ+vcoXduVNZzLsfxbuHez7DAbXqeXTT/LKxnRT+eDSiwXyk
J+vB/PZave4CPp5PhdaC/IZnIRhNpNPyH2qQi103HzT05K8hLnud8h5t005ddDondRhOY7Xy9o19
3QOeNg59lBvhrjUMehs4dVkowjVE48jY9DqI8iWbSa0f0gzql5V0MrLGx9KVm/CfAdLGCqBYVh2Z
5gHtcUtVoB30nB4dPH1fa7G7wyXT04XiBgJdOh23O5nYSFL6HR5sDOi+7zUfAEuzH9TDHhA1ETku
1/RZJwbsBo/rGxpcZmaJb5DY+dX1y1+JRcPceI8+ovx++BQhm+g8cDBEA2VDOQNXb1M25pK9NIsz
fjERirivSrx6iCsR0moBdsL1+VZixLErH8xipFRvncr1g20qYUbWhwTHHsdYBPExG8cfYbGKHWPo
qkHzIelByIQRGG/lw9H1qrv89l229FbRw4bMOfivgFvMa/5BskOEMrAWDbLOpGD7U6CX8y/J4CbH
2ilkjo5aB3pUqZ7pfMywN6s5vF0bFDWrrxfEiAPgzd52iOQ0L2ctEWde0XAcxM5DiHpq4n6Kf0cK
q+T0mfuG2s2BrQtfaLRjeuVxisw2niEDr/zPoCO4r+gfiF5OGptQny6DQ8bMjz9ZJAqLxpCYy+d2
BMK8Y4bMdvVB0FjhGGEX0+JPoySNCeHJZOgrU96wXdjqYF0PO/4qH7tO7k6oX8Yomqqig7q/boQh
BO0z6H/3i5pCKgbVNayd0EarEcL2R212w6at+g7QnTPnfnVgME9UM5kQv4mxiZ+uM4phZfYl1goQ
bhO4uiW+IrvInW4Gvmn7WmLFdMbco4+5kwoCg5NMazUm9vXzQRkBkIWzU5v16gpwywQBDz0CvQu2
nGz5fgm7OTliugKp1SPZ7OG1i6xvoC39NLttcbRh5usP3MnetC4yBf1KOkX6mir4ZDrVU/o7J+oo
3RF7vOTNC4FhBZRvUFXLxKYd2NEG9Tdl7xYopajmW9cecx8qy5qgPcBAPerT45XxRRj7MGfVLj0j
+FIoyUaLbXPvcal8sNGhk9lp+dJVpbDe7cua8vltmi5mxFCCyPWpq9DzCgVRc7JgICL+5IBb/XQf
1mi7fMr7Qq5bd6zWfKWQuxL67B7RO1oK8DvadGqljE3BdmqbNjsoGEVX4ZgGpPq0ALaHJSl0mwc7
w2lsx2AScSsxZPf3M/7jaFRxnPyOsi44rq3bxfcUqlwzVu6GQdBB+Wv2LoEyfoltKwbl8P7rOSeY
v/x1xHQ7QmCtgXipxp0KRtjejisOIWF+zNOYo7hjjcT9jZ+ImT21DIkMlfoig1gXfdUayZcamMFt
xmBdjOm6O0tWJqNMzDiNRcv57ohdb3rRCBaqYqoNMNk68stiPE6NWskmnbJRxYyaRrhPx5FVXGBQ
nE8KZ+cX0XpDs1pqSTBwhpXZxm6hYXz8iwOg/RpNzlttY0qkgIL4jY0/SUEucoidXgc9+B6gjvAz
4VCU0rN1BQvSICJPiK9OEszwXzurU07INjF3oyFfjIzpfcLHNLk9GTpIuP0jhVn6iI61rYkYOjAp
MfVZYYi9aHlfxXy1LUUVoqn8iJ7VTOfCOJ5cAFY/AbsdhchQTtpfR1uKzsamPwD9PK7Pjai+epoc
YGhHFOEDss3+Iyuwkg5blW1ADLyJW4/2TRWkKCXxkCQOZ6Y0Xsmxg4H9GdFG1KDer9Xo8wE5Sfqs
hZBNFN66NkpAYsERYvQsIVwhTZnIhKGzxZKlAyCBrDPP0tWOXHu9HSdESyHp4vHTmZSTaxoa3Bnq
X70jXXo9Lip8EMsu35yiRUqiS/8k39dZ/E9LA4RPEfdiobV7DdfWKwLpxkp32b+uhMyAE+LMQYK7
9qG+i0ztHdHUFBDVnyM1sF2oEHw/cgnw6YdYRQCzUHXiqaloUOZNGD4vYZUe7hqUdBVbAs9C4ILz
uOIafXY7sYLKk6GKCRvjhxE+Zwo0GTUJbYW6pWJK59JViLlW+KVfaHAbvDhuY24FtRjQUN8IjpCi
d6dcfhSMtiWEWN6DdcZMJYwmyBpU+n+1APPHOy0KmGDhR+3tlpA9StcJ3ib2Y8OuLNduXIf/GQKK
mTXfrRpYUBDQRaWlFLHUCQHuHi9nMrBEiJyFu9kd9zz+ASpk3NdhkE8VtXi1RMi23MMz9ud6nNp0
NChR/D0uStWiDWTDl69l+ta4y7VLlvdDsDKQuMdrQg1WrkN2yz1oJeu937Q125TtizWtP0X68ieA
2AUBLZERYY3TmNhOrHZOlL6o2MrdRi02f+jzfbFaG9dIr1WUW010T6pQINnmJpCvmhl3s/DzNxXJ
rUIxNcju9H4zv/CkVt+KzErW9dwqJzhKwirwN6NeG4p4JtpT8ay4Ahmfwq0Kz/4hXnqAZjgn7MAN
59pVan89C+SLAkiY/6u/rTLY47F2/ECsjQ0id2vWHRCyoIIKWW9rZc+zRPzIbrUv5ASGqd2sDQmK
e//J7aNxxZawmDsgpTRnaziDPzGOm3wncxOxV4ErO2Y76TJVJaHM191MII6LBuja9l4LHixVZ+mV
EbPb8661D5G0V0lPttC7hhsvuTyfS5/iWiL0OAnaP5R6Vs3yOYNpSxUHppJ3Vy58Gr7Ie+Kfyz3O
/pr1gtT0IizZj0BvVecVfxepEQ2eRr5hg214uTgn3nHcHBhf7q6JYQIj8Dvm2h/XzxD3vGG0If3O
r8s7anLJnBu4P6kc9bSLhOZpLeplEerLaUuUBySd0r6NeB5CpiUAgwGZELZWPyeiKD8iJWxA66pH
/X032CI//609J1nrboOy9zHe2YgUVAqzQKpalktFpmJoO8rW9yKh412+ZfNtRawzVhN+Esk7hHTY
0laRFUng8DyovSUKvEYkUoiSCO2MTa+m1ug7SXCMs8/K4XGWlWR+oWd9R7YNvA3ERNB4wYD0qzp9
tUfCjBZLQN61wBmLwjbk7TdlinRLZJkXin7mH76pLMXoEPz6jbOEg/7Z7+BTuFvimrQHAatFPg+Q
VGEs32DQ9WuLaK0l+29sqEhE3DyDt4vxnNMSZYD5PRiUPrPUrwuSkLFP3ZTEXWJbYfu0fUWvWoo2
u+jSoBMBvh3d2t6OXuZlW4Fdcbg6OxdKycvkziqe8njn3PEEFjoo2OXRUi4v8HYpa536w05u5uRI
illPwyvyxwFXKXf7eeSvIJDO/tvJdHe2QguQ4whXZ21R4ly/ABu8Bi0eIjHeMRVsRmKjMl8r/XKU
K4D66JJzWT0FL4dd4gR2Z3iSyGdR+WppAofhBd8C153eCJ1e8aphCddNWpv1Mnp5TzAu8FsDmSv7
zlqk8SMdepZ0qYCw1Np6zfSc4pmNdSEdPQUokc4E0di6t/D9oqiT8kdB9WBmKyHUIkx97G41OIHA
avzpqtqmezIstrz4l+ZiETT24E5X+R39rQIMoYErGEwDgLPFtxQvVf6fKzMZ1+x+LpX5Itsdj0Fr
PrFe7D/MsHqr1G8Amv3VdZrClhiggrf7T34CyByalj4n9s8rLW3YKt4VuA9sra8wN6UMc0Twej3S
VwvEwCtLOM6Vo+SGhJ639IEiDKEN1Q8sroYTyktZrJq4txbmj3+5M40Rj9fqk0Y60tRXBurLnGth
S6zcxqCUmMLPKo6x+d102c9w7Fmd6sC1rYFxIEFFb2tJuz88W+jjxQnBeOqj1vZNzRRdyU6HdIxg
rwxGOq0AEB4oIR+mOAtfCW76XjPnJoyA7hI89MY9WSYIBn/aGwwXM+i361jxGqMGOV31Spaeiukv
OyombEf7QYihjzQzmzeQxMdm4swRiIezkAn4ksQA3uBMmMwG5PJqLkcg5BU43sW5ji+NYMHJ6eQi
+3e/GzVVMA436djNNufLfFVEkKRIJbqRX7uMgCJrZO8buQ/rUxPC3oSdgZt7qDpI8/xL6czUmgC5
Xqg2O/ltbNTANCCc1uSqFngZBHx4xV/oXTvMCYqJMaG6PjW+MZJ6Y+myd42y8NW5s05bLeOBiO1H
lhrO/mQ+seRBSOj4JUsd3ysJFY/OeoL7JMDyoycYnHMC0Nz5Wn/Uljg3Ees/h+8OStDk1P7PMDPV
iEyHZykcvUEEscjzcEUCk+k/UkP5h1Btkqswr0/xakYlC6/i+5P13r2XfJADCwoYfWo7xrQSmCI2
YzijDoq7SV3m4nYp1o94k1HjNiUNsp4Iwn/6Vct7DH1WV7C3Fim+HU41CuldgTvPZEVm7AaLPlcJ
Z+iZzxBOvu+jcwfLencfWs7+ckVbo5xeKxhanQu/3pHxnS7H0TFr/Sfdf0JS1U6WfuhfgyBQmOvi
1nkNg8Ml9xQ5bhJz04TIWfdzPGJXAm25W6yDiMQhk6KNG0cIW4HPiQ+y50E7mutDYlpoKTmzS2kQ
oTNX+ZsyvezengYq1EAh5GkJLDxw7o6KF5HXirnvwLs95veQ5Dg6DiDfWACDN1JPsrHq+Yz8f+NG
4f8+8KMwYjin1q0bcuiX3Snc98UVUp8SYek4MKFjsjbXqRbObu/TEi6nJdO+ekdTIB2HD52RQnUh
xgu1FNUNQbnUW0MiSMW1b7gzpRNclLKT1635ZH25L49cd9Lmvb2+53AiptHyBxGLqbgw9xqFM4op
uaWafvcopEvoX7WOUE2JvVyI7QPzpLe6KpfJrkc2Mye6NgGCwG/nelFZ2Lwh6tJlGuqrGrg5QzS7
ok9nkMh89BoZksdpVzecFGVvEXz8blejB53+YlhJ78b894NSMBZhhzoXNpZGYEDjJcb0BOU5HST9
wmM4iavaSd/PpFWqYBr3gLoMgnj/YrFCA4MAmLzbNqIfH6IIKzGKB0uS7lZ/1tlTHJKRQa5F8qnm
v0x87cHiSBRxXRK4Bitl+mURopDDP/p6/0Um3i79nxcSiwUFD01F225ZqG6XmKtYzmWEN8LrUCFn
j4DM2BV1xrmYW7tMQzCgRs23A5323p6EaSi9i2wmcwq47KK42XQZtC/9TGKIFCYIaaIX33A0sQeu
Nl3Jd62JHv1Xka1iFZDgTh7haNefjrh7quQvIVjhEEthNMb3C81mS8ixrPfmHm+ZUgJ41BeGw+3N
rvWdflgE/me8aSARo5X2rPw36T2rZ3b+voxIls81x8NnRZph81dsj/D6QOqsrlah3uJkXnzWQJBR
fH2s0aOJiqQxrgnLaDnEK8Lzxm63ZDPQSWEJ3VMDuzKPSBAdyFo4yzsLGkiCNDgAS1KDK10if2gg
F+XrIen1ZpEysmYiGzji8fvQptCV3x3j7WFU/QHUFFSEZJgUgYaojcZsGojyUule+bbyFiNn2xEg
Ey4JS9ndLY8ZJg0nrZ7Q5LX73YIiYjbCE8S7uXrxstQ9Sb6BhWj1PDgv8Zt9ELk6abeA1XpsIWOq
l4zI1Q0xAGC3u7PDF6IZhQnVG8To4bRHoxq/JUNWXmyKa+IqF7pXNH1bWI3KmMIH/qOs1K70u7Q7
69tA6UXUwXLWAOkIC9ICli4x2GiWhkM2X7XZvt+Hvm1LlvOYu9ZbN4hrzOCOqlG0vMHE/PHIn49e
DbLusKQ1YYfsGq2cJUMnIaSaREYHwIGUeyZr2qB/1AOaT37TFAJt+QcN4/wM47tJybywyniiNplC
n3kktz492V13/8vylZjYQda9tUWgP8GXMg5QIMqAyJNfu22L+x4mCIsZo7bxxSARY+na9C2IGPoK
8AjO42laF+LRi88d7U3rwAcwu75KEtqbiweAQpODnZST7roLtbtUddu0VkMJzB7SoYESIj5DbwNz
hyZQteL6HMYRx7bdd6RXDEKcIZ1yUnngPyOisVIog6zgUbG/kaPzajfrYggWoVrZXBzWY/l4RKZd
e1P1lMx4R1j+pj38H+M/qbrgXIb8chIXklqkPSWv6tG2zjlgzBq90zkSXRRD3jA7pImCHEv+tkAF
o4T5Z3wMOg0T+ku0zkizNFzoD2B5KQ4QuIjupMUGijXXI1qRRoiwJSsDo3K9PJINsQdGKoT28tcx
1EtifIAF9vbJCq1BXbf2FYQTZ0RFnweZpUPVCPNZ+LKI+VoNLBmZ8PNB26bd38PO3zsvWC7l/q5d
TDxNrjJvCczOqIPHbc9Z+kij0eZxx06JiD8HOTB7sX0Ew04xz65TspVOEjOSzXHeL6sXwnHefQh0
xPI/PAZoDVuhtXbbMX8jFy9hkcgQrTkHTt2kfSfPHYmqbxeIs8h0uAK+PfyuXGdAV7XTryveq2Iu
MJseyKF+kdf4Fky3m1XqEQfqoc2RZUKBNKhrlHU1Pe1Ukn7ZTtV3zZB0dxUsYQpi8+nZAqhkRCsS
Doi0BSN+1gUUQk9N2qfU85OaBj51DfH8+r79NAc3EmPamOs4IRsloI21jLnBzHF3VAzROVwd30N8
neyzTXSP7xMyOQ8tNR+JKBisT9a6+LrJkpkyjVB03QWx/nzOZf+2Ahzn1s4kDU7X8PDLDq7zBLrd
mv20joD+aAxp38ZwUn+sug4+Trg44UtJvSYDfKwIx2vjdGraNN7422T12ceMFTN9JVJyKCvNc9BH
hv6qarFEIWPplq3tAfHP/MZjw7SPH4J7ybzI4q46VwqJXrKNU6y86oxsoOHccF4b/4vImFjtzDeZ
5CEXWy2BzBsxGRI38x1dtwmRChUuSyK7agnNZbOEemnlTDqWUD+1yLAxrfzBCLYcXuM98x3yZjvR
Lnxx1nzoGAbVXcZryPyiMTxjrBuUhv+mDFZDDRxJy+PSGx7scnkgk+LLR0HXYgWXfB6d3LSzksfQ
+a3CkIN28zFgI9zZ4jLTesKEdet1BRo8WCpSi6YZ3aItmQ9elZDfJKFrgHuyGwVCLwVjfnDENKpb
Ydys6Zt32LFncZyn8O9VWrWki8Vf0Pe3E5AVGUSXyqAie6U4jdY+DnV6hjbhlV4x8cksEjyJjwkp
rTS4W104XHJaK1eXL8QYI2Yh9woqjcuAWZG/Zyq+fNl+L7J8DSohrL5DZ1xszg2QuRo39i7Cy+ip
fl9UmV0d2ifqukdFoUjxBzsGUUv5JNVF0DIlBm8FpQ8EuHq+htz6bH6huyG4/iE10kRywnFWp9Bn
/XtOx+wjtDpLmH0YIgYjbAHGj5XzTX2YC8KsEVbXqxOrWrOf6C0TbPjvHx1Yvrx+8xm2BmR7B/jq
x5GJ34x+R0k1uF+Sg2dIzLo/awWvAPZ106/o4QBmON+n8s1X6naIf4uuuiF/TEoM6aLR7dtW7gE2
XwsN7OFl3UMC56F8PpbnlpqB8AyQ4jvrYff+kUfyhNXgqsUjTHQIYyYCfEQ4iBYEgHuPuDs6EQsk
W/AmfCBZQ3P29IjOM1ozXr7HChtVD10Yuu0XAdUJotf2H4Gx1wTLWPvS36z5FZhL+e6WNd4FpUkc
J7tTUXkA1jIj1gVPFQYoeqaVQR6+wNj3mur6CfLDSidiuaLF/xsWkDP9Vav+g7oCRB/Z3qquQtwN
V+eikA7E5fukMzM+W3fHbXnSSSdFnwWK3GISimi2BDsj4srvGY7rbRU4RYMvq9i3krm+m4hWy96c
8xzIigxhJJOJfjVVhcppqoSIKaHWxwFFSuSgE+Vy+w9gH2Im2SNDnCG2XtlMoYyG/kwHaF8qoggz
RmIA43H/n5eoHRYf9czueetaJ3bvDnqIYmMv0gjz5hcxUFLJdGzt+V0lE+ZHC1ImLAX8VFRQfOYn
1VL9IsajdU3JAEw45gaH7LYWCTHvj0Dwg64gCdtsGIsY5J7tWTwlJhxs+JuC1axvWhBElXvw2Crd
hErpT2AAVItT+W93L+8eCWMRaIPTgQfxRMrmOSDS6oD1XqbyPwPCZzL9kDg+LkBjHzrXN1pgCFqb
rq5F05HzU+uViHr1mFONWoiP/JO4bgbGoN5wJAyvL820yXqYg60G6VH6RZb/AL14/gQafddczpJb
FKsNGnu5i2tpe41rQsqDY6bu2K5srXq2BX96Qu5LWBOJYY7e8yqEowldZ645AhLsrY9BD/3bosKi
/exL72FqLvS0kBKcPWTJH8img2hhKnPxikPJl4RNUG3rgUTNbW6hee2u1rgf90F2IWABw7yBCPqL
Z94h92h1/wcA5XO+5bgFkUSQApmiUavTUbznBDlLj+RbsVMjvUOqXK6/gB9TTjy/s2q6CNH+y5ct
WOuwCdZQvFE6cDrUiGJUapxS5NGolG+dnTADQd5yIgMVMx+TbTk0txpmo4AEu5cva7MTqmxl4Cex
J6JcwGWGxiwymIoeggAHo6fzKSd1Ui3o8kxCucKns7gPFj8LKvGjR2+qlwl6oIU+gy4u5drSgnaM
WC54im/2+riVQm4lq04HoS7DG2Fs4hpKlgsEs6QqLqKjDxZXL8Bvn6rgriwl8RMBk2vnRrhPc1xC
pJo3XQGS6I6CyPc2GWuDdvfWlECYGtaUlEggbfQjhSHOKCfEL6XZQGlSAcpiGAqi3zRlXt0dcXzG
MKLeQUyLbUBUJr/9VbhaViaIr+ZcoPqSiXQOX1+vQxk4yv506G+SmfTPe9CNw6UBxTzYIajJQoG5
uI8gOgsQKWAAJfMQ3bLYmRte9pCkjLHPkBECHrbDcWteTe4lY8eY6hZVi26xaGf+nAiyBBGsKPpc
E3O4kLmysyL5ZUr1IVWHxL+chMrvv0TiYxW3/ORL0BVr20Y+8wExXiVrOxomodi0RWXDiryMMUyh
5P8Z2MoVUzPmMyg+z/BsYAJvUO7MsH/2somOIMSrZxCSj/G8IsM2DPmAiak4B1RN3C7+EjIj4Mdh
27hm+nhc2bt6b/5qLesGxxaVse9LSS+P0wLmVFKlM0vNnm+V9BHAwfGhlEiyLtZJN3Q+OU842ZdR
MeNMm+kuqBm4tlWrMrRA/jHkckQD+GXh30h4loXC2D7btQO/qe4zpFQsUzcn6ZI+AJNLnSjI1QpB
50cNATkZKC4kBj61m8HRCiA1n4EGjgZIb68yQWLDkTTi7SpZ+YBxxmS1CR5Fiuofv8WBBcUFNKiZ
y5j9nOaCoHImoTR9tIdCvI0fUWP5NobCGbBET11j2hd5u8f0R0MLerodWU/Q1485fVoSygKJEG7Z
wDEExKSqi9AsqkRNVj4heVaUBHwo2zt6S7UwJIhf6mw7CZofwRnijcth+G+gfI4RM39TNI8NGZ2H
zVL+w1ETT7Vpfu+klwEh0CEcEiHd60GMjhDNrc85Z2SNAaxAXKaxoRaZuR0iK1145BqEGKeJsS48
2/hP5GY6K1IW1y2VX2vZqVZbRkNLDHGlX+ZcCQ0XO7OhElNSreGcpJ1aF2B1L3en2+GtlyS1/jS3
yxH92PDfQ3k3UJLtDMPzWTReifmIkGW9FGWTnVeDRdy0UGKjun40fXWxj2O0AU1yb0THRT0aU+CL
D08IeLAhfnP/fKOqgt3XKBY8lWCUFSPfrDpQWR9tcSV+5i1oGGSDdBF7Fv4Npua2+eYKrsHR/qJA
v+MOBUrIRpQ6p9e1xZMkSDPXpUA4OBnVkYmyiZxt1QbyyVdffYGbDiZpecCXdUENMK1JB8PtqRg7
KLPKybmGAo2qgKORuXIdLvP7B3Mf0jOblMoQqnCjXIEvrKszIMUQAa5s3FuncAoyhM9rJv5qqCAX
2D7F108LjxneyDkP6H5wxhQ9cIlJJOlO3pm0LMiPvmiqnMjoQtYy9ZQIhz51AAyJILejCZfDDqeO
iQXGXsnBU/8CBde0l+71EM2J+hZJTMMtFI/A6NyI9vByZW6M6gs6RSxgQLRe8oRgVCtu3nk/mC6M
1nBHBAQ8yAKuDNBdwGmt0xVUCfmb+UedQZ5PknMolq/vQWtBrMaVDLalywpDoBQpJkz43oQcehPg
RhzokiSbHL0DfI4pZDSb1nx53XXgEQghiG68OMabW042fg+N3wyEvK/ODvg1KK8HhFC34oybR9AQ
o886FtjZphAkjwZZjRbfsoE57udqWlpyLfNRC74HE5Ka77U9f2U+iOB862VTEa1JYI+TxYw8JC06
uCo2dyXIX6K8tNZT1nCAGixjBATKNvP130kSSku5n56Znr62SB2FKfycuMa+FtZStL1c/DhOTHle
I1X+qLYgpyhmBhv5whXVtS9YZ+IC/WLxgoq2sjaE7bm1M+yNQs1wKpqxmaTziu7LFRvMtiO0tCq9
muIyfCsMNqIlcDbNZyTr56cRr54fp2RXv/QNR3uTfkeNoX47Pf69fX3dog+pqgAjfZncGHOZU3ql
y7ujLiTmmOK/yQQmIOj4ydpcFvQOIfDkEgu75pnVJi+jE1xCmAy66kY8i3HyjsxgCBqrvgUoYqJe
k7e9qH9LxmGEbA8AIwNU2ScQW65RTxqOcP5zoA5RiAX5U0AMLH5Y68st8ktn11qV+Au4gtncUWtY
vE108Lo0Vzr1Ny4CyWLEEaGwwlZeh5Tg+/UYcW2KVOUtd+NBIoQgSDmUvsWwCI4J/nQw6t9N8CQ3
JPEf3h7AjNlZhbXA6qB54LQfm+5Ml9/LU/rOByAtN9qDAXnvzFD/MkCWnoJR2OZHaGnwA5mQzo1F
lnNK2HeG/OUuz6Hx9MbFQi5hpzGEjYn2ct5B13GJ017WFO1ntTpQsIyoz7UFpGNMZY+4Tx/7ElBi
v1eN7euelo31Vy5TUJqUATCR9B2hgZvB7XaPJSk9LRPs7WtO8yBScOe+fj+sDCMj3FE3++Dd+1+Q
OU9PHPTUbwe/CUAurzpifGx6DQKubN899qvjfhUVkkQ65dTfXD2lIQ6i0JrCjX3CyE7HazMGm3BW
oG9wJyGtRUyws6AI8Ja3DR/owon6q+Xf/qbL2TmTB9INPD688rwplCYIMw0N74QC+wXkKPcqwchJ
LdfqCMvkhf8JlWqB/P4RJJPtkjsxIOWe0oWlVNF6CK4ZhWXDy2LJZnlllxJ8n47syu75AgSw2tCR
jVhWyMgEBRIr4ILd5ztHvUg7iqB/E7ILzeVoGfJryGeUDdDBwia2Q4H9BHK3FH+CtSDhiAw9rzYd
JapFNpiXYRzdl7tQuzvJv8cKaQIxY2EL0EEX7ASRIjfkByf74lkG8jKifbWc4ofsZJmcSYR6vI6C
AoGqa9eIuhYJXpgcL74UFFlPnJ8B4Ac26Zo1lP3+rE+hBvulAKVYJEyQ31IjuY0ozepc11Sj/w4z
DMuY3R7FVecRh69stEL3QnDXS+VQpihAondKVzlQyI0kxWnsi9XwjQnI5KmghrKB265yzugwcjXQ
pkLUpQldSZLXmoy8o3sVOvV1rhMT8jFVaMRT1SjaTgEF8z7mOdrBtdeauVpxkxR5t6e9J2bGvVsa
M5d216PKRNBBewOr2i6fikDP4BFKYtgnmVdacWkxx5M/ZO1FnKEIg5ulWtZYrar9vOJI8WVZDKZv
iUt2vp1ndSO7Qeb9Zqp793idBCqUGRPnWZ7lmCNmT8o9tCIQZbvM+68cWieioqtpImz3Sb4tfCle
stI4MtQYTg+J+wgqb8Ca3ZXcFaD6fQWSWkbq1hTWD+U/Ig+i8sNqh+Y7oMvPKVsyn/9UdDRX1B1q
lwyEgYCYsRHZVXYdVwH3iRHSp8ro7Cgb1p2OkQ7kjmhU2sa4nrnlIRJZxF5QsvAQdyQafF4adf9I
Cxy3PPyux6FA/93WhRj280c+VoW8xhrHn8SAw/6e+6bJxDwgpp6mIhhQvIRzXH3LnWbsaIHOUUsa
jHLQ3f8k+xBNokhHPljnuiz2qF3/QMzrknTgokpNmThv8vubZLRKMFTus837TIL/8faZcsqXZnBP
4NOYE6/KwbzwvXZj5rrIYd2BbIjr0nwacMvELd9SVjDxogu936gUmC55/NA1xcUPvDXllpoRpOzK
JzDCeU2C8Jn39zFn+eX5efJC/skIwasnkVcERK+NVBObZX4InMxJcP/3PxVQUKZ77yym3jCexUuP
JmmhGelIccCVrdG+A6cCbba8P/TrV81Qj83Qpl+arQhhCrAZy4VFv1KA5ZZSOTqaLvmzVzzMa1kl
81Gxb6xaw1afLBNbci8b2qwNBx+8uct6O5XdN4BmGbj1MCnqI8/Csr3mHJcMaYBDBYplFEYwXRzt
SSEQ+jH8WtKnP3Atm9R3uPoM2TkJx9X6PNexqwPxNDvI/rwakDuCO1YynM8qCwVoeMsixRnyglaQ
p3jriYb7vc54kV28JCW9VQeN0mw+MuYF1NFIuJwfqoGOzgoNWzEiRL8ghmxBQUFMqI6pmdZ8Bw95
EJBGiLbUW6g2XORDmC9Mggp5oep/d58ThjKB3+ET60v7/NkfbXMGVTl5zmlUrcmuPAoPJ0buf9Ek
qDYPq4zTdvBZXft+WSfbcAg+newC36yTdSqj9aHl79BhH86q1JYePoSo3lgUPy614VYjlZs6jmLv
iNzQZbAb6EpdjNVOKfzdX8mWyxeq86O2KwMmy7VgL0ZE/d6YWnEJxW89w51Ca6AKyztr6erNGd1l
uuQ49+zPLAcYXsC4gJn6I1TLf4uRCRVIdDzFNuMXKI61m04eeAWnISAnrPRWpXDXjJWbn6OGOiNU
KBFqb5QbMyhdSI+a2XVmt3KQj9aCfSxr5DYEr/Uisi9u68EraHdlvQO5cAJMGOylE7CQ1SgFBvtb
sOSFDemUFuSQGRBzLk3a6ggmsoCWP4iOiBE6jE1anSGlycZS46AguPX7BB5NzDtoE4cd2dqueLOz
FvgBK+20hHSDoeJY1/FGDfgVVQwPIpy4M/GP5SsB8NluLSHK97ozGEv65jvnhUNZefuHGh1kNl7T
Rrgk8vYJXKox5TsIVrzom/SyGl7AYRmKo54K3SymsdiLSWzinhBMCmNIV95q/xaKYYQT0/cuBCSa
hrcHJmexr6wBzqoxmpFQ9Cg3ooXRw+1z2qDo3BQVEy9a6FWgy+sxxEQF99+eg54JdEYZiog14+W+
27EXayBbFfGPVpBK4Q/+eJYOJ1JQ2+WQkoKftbYUiN3J9JsyMUX9FzqpJh29JGIMivItbZPjak3H
/mTNcBvP2vdyKXqhjIpcUVRRA+afElc4CiiKooXVSfsSSqjAfUwelq0Vsn9m5mBeLF1siw/lGMkh
19VNTsNlz0jeIPazwm5iHLm8yOyDV1S7e3T0018EF62OA3Uk+LMHXltirLTFgjPZtTj/VoshVkKD
iW5hQHk8+6FUnIR7ugHC99VcHHD5t/heLk8ZPfXB44kuOw2IsihDPglTYNWUn5xjdizVDC4SRwe/
cORtncjk5jYa2I/pHZrhHiCGo0pJ+R7YrKmsXs1YA7CqtTk/Gsslmz7ho7L5ZSf1YwmjP7mK+7ma
S17rax4bRIzemOX6BBe2x41NZ17Cemos0mqwilbHqN2ny8rOqUZo2IOjAUJYAoMxLo1U7zp7uQB3
ou1G+qp0XtsF/qU2ZuZuzYkoyFAMxM2Wjkxez3yI0vDzHobAL1qra9HhO2EYzJ3lIzuTJLrOKqFs
DTYiQM1G3V3RgSZ+q+u0aLuarJxe/GXxMihpyOXd84kVnT838gs1fAkHrMCb0wac0QfR0hutAAqF
+ySkogJyhJt7b9dZBr70krP32gtjiEDU+vgUBKHvnqRfQkQV4a1mzIgjPP1TdlvmHVNW6z/VztTx
2uJkSz+EnBp8FVB4Y4oGi+WcAQRrPKy9P7EW1Onh/YlltkWgaYifBH4X/Mi16InKXnNu/zUZsNtb
FXb/GdhVasFL501yQSvXM9WcatyBrghHF0QReW10xNOQtk/cHdcqjaDvQMskl0o6HNRe9/cwK0G+
yolte3KZtyZSSe4GGRs59OjxFDZD9ewDzojJB1zx12z/d5ItYU3DjaHJHgnR+gVEZvShhSPBgDAO
vDIPHwMDUzVbRHsA0/q+1OHqzrRgzEpHM+BkQHz9/eBV+rAE4DEFfdaETgqAY48PU57tZQGJaTqJ
qTog6fOsn0rg86oIxpEeEqlwHoy19DRmZ2SqghFoA4XcKvXUyVbg/O77jWhn1HkeafU7JlDsaC2k
OZfTX+LfuGhwuR37LsgSsYzisjsST8FS5aDRyhpyPfaK0FntHrXtITT+jy7CBJT+Tsjd1kSqkqbK
1i+cSaQCidTk/+lRcZgkvFNLFAzPwQDeRBW/7AFoTw9TntlxxiXjKWp2RnS9IMvbCSAB32lm/ryb
5feU16w72W4vN8sw7UYaIUPxqYbvwpm6Nn8/kO3HVjlYvIcdEMjnW5LVErAzmofuEVjfjnQa3mvO
3Md3Wu0XUc55G9a3Y43xCRjx73kZKklWLZmEDvwjiTwGYWsvDNhgVq/I8dQUTOSHnovGyhEUjFQT
JTiwPPPwYeYf9i6qIS8iLkqHRLZ4T+WZFi98W0jIMDMIhzpTwtItZnPV2NYnbEI3loKd53jcnOsK
YQJvDu+N4M3bBEoEBrGI3ygHuVuwee/VyBgoPpEB7la3kslGE6aROaAWiOvDiS1hQCss/4FNj5AU
4PBfWxhSuirMayFbFgDEYLB555USvXjDA1QTA4xPxoaBURE2rLvV2DjeKBKLYuK63mrwdij9nFjb
ljamZB+byeX1mqhSXx/MDLB2KWgHMzHUjsizHSq7dChm7EA5t0bNYMz6Z3pE8fk5q2V0vsNfp9ag
By7yNi4BhTplKTlas/O3RwAbSTbg+HL4aL3qXgi0GSt7FT+Ig5mHP4CapowBFLvp5W+JaGSAOVco
EKqODQwa62Dk6NL9UeWQzZcgOyxI/h88N+MalN8uBKvZ2+a31XF701eDnxu9NiVhEFB8/NlddCop
lInzN6OaGRFyDC62hGzSBwr3kwb83j1rHNWrG7pB3QMThXkQoLes0kSEdQUgd9ALtv1GrBagl4TH
3gBuCOXkskWjdRTjzmtSdw7RV2cw5XTG3Z7MA/CjqXMCPmaacyQKoCbwRMsFYieWoGqGfUGT0As7
zJmdKCXG/erJZPTWwXA7Hb0bROhGcC0KXa+Mv1r7p/KG5vB2HJvfnu+ws0ch0omnC5+Z+CbI3vdC
7ahvng794qDHVn5HdIdHV08B0tLmbdwlJXixZIw8n2Fmk407LuhTzxwnXTWhSM5DN63cU9uR89NH
CrvjD0t8D6LBYAaRrJ8Mn7bdnAV+1p3pd3BguPAitaEftroPK7kfnTsJlEDETJ8BYnWHuTpJrx+X
Qu+yfM3vY2p0Xc7FOmPxo+c2ZwUErLMT6QnT5di+nQG2zbzvrZxsp8KYL+AB3b18h6ME5vytALYE
lZISsI9Qg7fHZHAC+l3JNuVqC9HLVXNIrQ+vr1LeemMUg5ver8sOxW95EuD6BZI4yW+GaW0cB9Iy
9xyXidHKxlkIGPEPCAj0kkvxQMkKAo/BgnJeomlBJCqYsQ2Reniz6lsU31o5vGuOGMIRgDC4L0sU
mc292Rs5jPeNFuv89DfiQ3gsIL/Jw56pKnhMY7HGKM/mr9QbWKRylez2rnInBeWFRH+n+NgaSgID
jeK8i8mLuIjQLG1v+lIECBvwgQGlzTee+SGWStIW2o8jSHaMxIEijlS0G4HnKZR2amBhBzJer26o
4oNUAhmQRXyQxU7wx2Pd1/31DxQFF0ox4xSD/h9/AxWyLBaC5sg1rgApKG1m6L/jahRfrlIfeQvb
iAXIvUzFNsENfpjuw6Zd6KD8zwJNavP+WMNm4tNbmwuIampTSxuAicEndhP+mej9Bd2R+wM4CjK+
0p1jtBGEQ+RRGHHBzNnOSwJaOp6HPgm4SVhPSvowJHt6NQR+8aRCWZILS1rDmpQ7LKRet+fVUDvd
QwNOm7CUtl6++2Uawtwkz5sMUcNa51OPKP43PzFrxa+SJEcue3P6QrXzMk1VAYxH8UGpgevQa64q
9+Jtg5lhCeYO5heSh3eNaDos0KHxKucIfH02Wl9HQM65mBhbC9mZIu+pSPlkGZhkHnsu0uuWSmyV
p1WZmDUhzoV2AVgnznQcMSv9Yo1iXcpI7uPQEKCcwwEHc6MONWrtyJ1dp9pUrKC6FCbC/i+NcL0J
i0tGqIjofDfaf2ykQXx67cdVxR0fXrPRUE52h8s/DejkVGqHw54O1MR5fkazStr6Hg8aCTZSKcJg
t3IPjIdu2Gtx63I8FoPdxrshoYVgn4mPlqypNW2qOLFUeDjxHSVMQqvZ32v070axko+g5VeRSOtU
LeIzd9P2tqfoIaaI0XJsCF71RZxwd0Ja9KDnrM4qqjdEt0D4KQFVAvV1dHzC8MzS2eX/c0pAmIT5
icfZetX/CkaqziNqqVxPxs5F8ykuNjifIW8skN619Sk/yY9EB1+RyuI/d9GZIfi3GToePe9AtdfP
7tQLz2F3I3BAegLMRy/8DJTenCdIvpueiH80HQh7ahV61DoydMtlbDd/3kkBVLkly7qJ2FCITuRx
1iRb67s5z1cioSG8tbe5+/HSL+/OHzLnwyUjrcAnC/uosx6cTMWLdB+yCNI8N26dIlz1afOp6yiS
jSF4/zQtYync6WW6lhWkwwBzjy82n3U+CXinfEN+Kmbjgg9N4cdeg74lqnuEgpqhGTPS/WMMe8Jd
AeQFEFnUidSRUV/p/RwQIRAVM/h3ZRc8N5FbUBTq9C46eBQ+s6zAvg6kM40mC81030jpbX+JavtQ
SK395Ms38LlIBVs902GuK7NOLh77E0kJEhU3vN6z+Rzge3N++cuiPJvIxZZ7xNrLlDZfDNzoRVjY
wui7WQgSx6wbg4bn+LlGVlthXrufvofkQmk8eCLzIdlfL6uQypO6mpRYFN2C/zPuIoa59RdMgLd9
yvr+ObuZ557CBSrn1IQix/p7iCpE9IjwSvoaCdzNnbxnCgUT/fqQZ8TuSuODJtNpb4FH1uLcf2wq
CEsmUPOfFu8qEpbpED9Le0+xLGSSXTkurLxfNPctu2zwLWfYm5QdTxVdiEk8inAGYlD9BtK94BAo
kP8/PDuIvBVFbo7QhcMljtqyBJS/PXNpPa8EBYVtGXFrlR7NRJJEv5asWfHJtIQQBZo1U0KVT6fp
5WlfG6ez3eoO05hLW4gNbDk9tmpQtW7cd1Croqy0vEDRAhuygGbUQFbjbCZZSUqNu3FHo4xZuSCI
6hvIOxhJoEXXWtFvQGBWShb7ca+ABbyORDuQmziLCL/dsLYocdGoFjGI9bbuKjvpcdL4Eni7JvA4
4uoyml+ffTUriyTAFEAypdXdrpHHTXUUgucqMM414JYa653zQkwG7LvHohZrmmNjjnrv9BYoTvrU
BtJ9mJXnbU2ReJ6nRqOyRqKTpwCX/faTrXwVgRrj3ZmE/YBAAVueU/6sg5CeDZLiDBUqnv0F403B
uC9IUxv9YufFs0de77B1e4P9Wg1x80i2EG+DxMF93OvRK3zp7sVE9WHMrv1xIW0aXnBMDJ3piUwb
mRHAI2cSnXiMp0SUyC5fpkX/ex7nyKc6FhYfujFoQ2JFsgRetPYkSe+AxlEvoTK8DfFE9LV6K0Xg
0rFsyCEiwHE//g98NVKHAP92UveJUhEkqqCUCniH2NN/qYBYMaj6KxjeIDy2EpI46zlh9RnLujFR
XiPs/OYxEjp7eLoAtWHLaAap3r6TW1/lXbxzMxTvi0XB7S2F4iXpkvrH7rtWE+e2EQ38KNN6a4QQ
Q6uZuDzZSpeQTOuq7SY2AnGfPegP7FeqXl9s0M6Mn4orb2nbk36p8jThlWxWKc3nvnFhoIsOHlg8
94tbY0ogLVP1zZSIRbBX+GYP3cPGOuUX9w+VA+420EZXQu37BO6YG123oc/2ySr8KXQnbi+ZqHIr
XL9Snw6KXFhcgO0iC98dg0QJJxd1b8ILsHzFRfcpdMAoqLVGYNO93liMaeDcUegItoOGdNiSvNu3
xB2otgZIMMaTBWPVjdwM8/qPbg7XOD72oDz580vL9hCCqWWaFNUOQxoQgF1W4FM4gLmHGstOatbT
IZUaeSXfN+Q/jfA/68viiHUPA1utDL3QlWtRt6DZ98c7dmNZru7Oi/C/0AyGD3Lp/JTE5XiGk3QZ
jcix46eIPtMOpL4MENz/R5lA4x9FuDLuvOo9Kos8KIz4mKp0fDCAwoqdtfCioIBB5seRyloHJ0dw
SNmHyU2CTN2qbTv7DE8tHgfp0AlPHHWsz7Lb9H33RRVmOUhPZSR/HG3lVYzmq6lUpG5vK+72PENo
X1085mVsbujZQAowakvg8Isuog7t5/xzHG1HcLG4m8ouq22czcJyCS0c31oZO3EUI5YkhT6tMsuW
TdDmNgBFyYDsBfP0eYbj4B46dLk1rmAuR2yhrBK4Luz1zz/3b/n4PG3aWW8fB0OBoJ1xDZ2b+bCJ
hDCUYxrMWzpamVmfpAdexqNaBDGJnlMUNeWnGBf2r5iAouzYqo4Y1pAna5b9lNq3pONSfog8A0we
YSzcAGXd4f7XMRoiZTnwkjTi0xklUWKa8Xq1vDdQNsZ9B+HLWjARR7Idk7VXLzchD6B5MMVSfScC
GkOqfArRT+YsFcYjXAO38yDXzlHGKZD2AoUDpiyA/8Dw4lZVi6KrqczU5VygJ15fBVEiLdIjF/Fy
pTTsvE1Qcls/gUHLVoaCshhkwyC6blouWlGQ/PntYCk/tDFh+VRkUDzwNbEF9Y2qlpYlabkVKHud
X6wkXI6tpQOo382GGhwh2dr5Dd/CzC8ak9vii53GMO/SKr4NvrDYNcKQYGkw1UHLoHCq3R9PpeTE
VOvnqvSe8GbiVMfJDpkinLpBoeAWpUp1mEOUr0Jq0FcXWMAWUwKkmFBlhnFI3wrwXTb3xU6Xmt7+
IocpbZ5yOBdTlmnr/0fhMjEvwenOhy1iTlNtn0lDmzYvd47OaAAdWPJJaizU7EoQAiEgYmRjV/vs
Aa/fp3MNE5LEr0vPbBK0M+ecBLz2xUiXK8U/EH0N5Hqg/c0N4G8f014LhoccbI6FcXZdeiXHReN3
Kn39ArtDEZqgOwc57vQE2srIpeMq8/DjHUQ2YO34uC3xYH+jzDtPeIkmzYgaMpF+O2T3EBEAM7Xa
XDN4+1xVC7/ZmtByCIWARl5CEufwP8FO6lElVuUGilZNtXsikbOryWDPyvcf7qPSID+aJbsrabFU
P9ojDjLeyNYiaCrGklceqqlPdBDCxWWj6cq4kwpQao7cmq8d0mflp07uapCL9LwtYPQarsRZIwTX
b+ZpMEKg85WuaxQeHvji68eW+K2qJm9FjFey3efc3Ge40tA8/++CRLeTJmBIR1TxMYWKhUUl4gEz
cW7mZBQ966xdNF8fNIi0Pye5s6WBYRlr1mEe9ocVyeFzSIVaDna1F22CGlB23CwUQF8K+GFIljcn
hMjVSZwaTSYqk3AVB69WAROhlB2XJ8UupyewZKwZYY96AKfeiXMTkOg3MRcYwGapOpDpC/WQAvvO
esduugCtu0v8eTpHtPYP7pnjSujsQ0iHMAkBKEaLv6HjS1fqzUSYrAKqhBVkWiIwViYn/rq06CpU
IKHC7Z+eG5VWfnRmxJLkIeDQTPfo8Owuy8cuE+WKURn/VsBQUfLymQB1e1xYjsR0yAIUPgAT5gS6
/PTRi6T2AE7RoiHZVJJKlIB2KErc4RXWLuDUz1BSL+QOPe8ve4b4zwnTurCcRDnJMbXyJgLdKLI6
e1ZZ+tgXQu1l7Is+ObbESdKv5m4pABYmhi3Vu+4gooe0D6sJuKi7EFD8fyvpCOAc+tRKrh/7p+GT
nUbn2ilNHHJ1DcgoHC5Fzb83jy1cxZ4VcbIz6mxhOgxSHsJi+eDiQktvSolnG+nhy46KbESsEfbH
q812lBnS3bEuVF7+V8ZC7sxXF1BxIi2wXPYLBrWIyOC0u42APVH++pgoum22Zg5XAzSSjX92Nq/U
4HvssDEkq/y2J5E3EgbSpKa8YjMAeHPqaW+OkLUKwWtKutQVWKDEpdEl4Kyrr0Yhm7j/AuZ7/vGy
CrG7pnko2yXByX6gz5KZbgdy7SEaDgyovCAgo9tXzPhuZmhI8OPBHpc/wqAYbBj4fveSFqwRR+Eh
C/rmDjtg5pvz3XXhTqjixxU+s+CH8FpiRCjIzHkGFXHxoECG6B7AZGO2EC1eWwo856/rXZn3SKTJ
owYLoyptFur2vMQpvcd76wz38wjRU+Vu/2QieANQAOrgZHPNmAzZPHXSk0UTCdZ4S3c5so1vTzqH
shHpRGfGfpnJKgA37aZ8Q7fycERWbpsgsdQOrp5cns0OxjkjYR7WwHb4F+S4nii9PzPxOq465hRt
ZVQR5ZLcI7TX+LO7fO5wzFBHUIIu9boPo4R2dxptkzzyQvMSA883MQy6riXMPpao2ePtmbk07pN/
mTk3vddyPJoW+EIS1nVFZH4K45vA1Hky7Qlo39i6k5aLZKKqggJEbPb3JWFRCQXX4OYd23rlvjcD
/uVSojVEq0v5rCd69Z1Dn+NzHL/aBUHZxKuloDzARbT9XoJT2TP1vzpuueopIp8i2j1DVtBqu5Na
pwtgyX660XVraHbt45JFl12q8GwMpAVK0pJDkf7KR460aNfa/nEqeD8xjRZa3eKiQAwsQ1ntPQwI
NMLduSqIxe6dfVjb15siMbknneCFpd5TTHNR0XLmMm3STfvkf8XisFxM/IHPbyyvrLrnppF1lEY8
zvRxZ7OA3SGPKD44DUe0KOUtl46TQbIH/XaW7bEcluAQozMRz41VDnNQQAM+WKswhqACwzECZaUh
C4TyEzVxI+28CEmGrl2v6m5W1EKW1r1wFCrr8byNk3L90q5rDIDsasVHs41OsOVCgFix4Eg/9MKP
0m9vDDPX1sjdjFClNVXsgifQdvcq0alz386vwt+g///tIhBho+BMovomGFrqH8hMqp2f6THxug0N
1C9Q/vyx1M02pM58Cwcvg8Zklsg9jmpD8BokBwi/ojcchFJOUj5JomuYB1tHUgvcnI5xxN+HTH68
NfLyXnC89SNAHIMCCfPzajc0+4CSQBfAQZ8atp02lTWs0PI5/rtdUm/hirltzAUltFOgMizfWbJy
vRoRTVAoOXhy/+OG/mCbLYHpX3lpbIApaMhmtYBeNqNEbEuNeQdRpXbphepvuy76Gq9SKv2j0yrR
QWih4XIm/Yux95z2ZecrcRmT+CFwuJXLGzw1lflG3RLr53yrx21oMvcGlyHd6uUktPFYZNoxTMlZ
d5JO7rH/IcCTivVBuRYcKL6qJrIlpIC7+LbtB/nLaNzkZHOrsRPJkCx0jUMjtEYRv3DwITVUPPRH
FJtiPAhk5bu4rpvt9VKQ/usUSJa0mhrsEewYyi+nnHbneVH4QRbuZXesOcFUncSouv/OZLOvEGRP
813b/Cx/ianw83iGF8dtz0F5RmuXcfbisrI0dNG944ZgWWeQeeb0a35sodyluR9CIs33p8WBuwmp
oTmQm4M64jEeQEKt0HTikRzpd0BGuHbH2JNhkKy8n3Jc4QW+SW7HF3NApbbASucjq5W37urOwtdH
ua1+07ZRkW+QIBs2DaJXqqND/CoWXTVhrISnrU9xjuAxt8F0qtTCYG4uSe+P6c5LmRmyGCH7/7ho
9BhMxzwMOZyd+M+wfaoOmELxc5ZzJuVvq2zQbC1TBYjwXUfQPqHOGJvlEXSI33xDkAqw/lvWdWpw
AbKdy+cU0NLzyqfkmrXL9mfWTiKHiUG8Asc/DDzRM7jSGz6ApUXFgVLtieBFgm0DMOxQXK3Tn83L
nSEefDDDcJeQp7T2tYIzgTMIEEoqg4yMCw1W73f0TOtur1chN1MdafazIveIKiwJueBXWcqoWNtE
p3bX3LCU5+jFahPezyv5IgTXF2O1KRTXdridsT3PT5SikOSJNbOhfWJWqWWpF3zi7XYs0tgN4L8E
R6/wptvl++T9DNGLj+sYrHNht9yPEIKNDrXB/aR7/bIL8mPZGphbCQtd/dpfYHVqq8HrgUvao9t+
gF/dsctBApv4dHVjw8Z3ACtkHwxvmUX5KAqWd3DKpKtvhK/jWLl4LUFwJRmkAFG6SfkAnE6TsTxK
bpGOZCdpT8S5GbuvUfTWyLiZoTocDu5y1V2xvNGMpGPnb19cKrHdBjK14bS8a8LB4bpom1ia9IRF
Gxh0Xt3yM5+wdQL6wa3FH27huNKahXjOcKN99XJ/lMgZzk/1K9PgmORWEx0OkLI9D/EFRn/eJIOZ
RQrsIwe1dHADQE9PxCQaTcdLpRjOkcVx85D4U6sQ0G5oYMoT5xfzdPGTDFNtHcsTyirg29ydBKw5
GfWr8PCBKVZyTbo5hW0eZgPykrIAj1MfVsJxzqIUOpbDAVIYTHEKFbZWd6Xfln0hOAOErChFh7UN
sLXYrt7SYMI/tg3hBo9PcKt0kn21eeEiOpirHf+UhB4V6o6NXdSJyCdvSjKTAUn0TdhtyQPL4pBH
paDu5k44WM+jRQKH8AVn+2z+0Uu1pMRV7XYKNNnmNBJw7BgrETSL/B3WHuMDehGln3mBaCKzR783
5mb850QFR64MzAk0vpzSfloaNbZGXKMmQuzP1j/Uh4fCPu+oS5lbVzM9HfIEPL1I1Y1ciB/zFjuI
+M07IHnLoKcasDvTK5VOVpp5Bg6Zd+DCWqfB7uoZImckBiIX45zdPW0Fh0hrALLgF4U8OcUpMbW2
KrvR6vHIh4tJ5DAeGaG1YSa/32KvVbjSTQ7ZjmzEiaxu7NtbXRypn8kHzOAM6XXq7Q6zyUV10J4O
UVxFvtIMrGV5hqak2y1aWtJymAN/QyMmE5XapMlmWoGWRGLela/PhIDV3YWRU2cNAsWKIDBYatfJ
ANwU6WDPlGfaBFojb9baITwyzMiZcDiM0yVZkw1DD72pRuC0MgjFE/NlAcu4HMQACv1soospGuCp
QStgQcqF7W67mw1NXfmfvEhKYFFqJ/kEIp2+JN7qsPcmaQWUl/lc87JK/c1ORRivcVBMlE++Q0K8
9kPhoQH0kbadsXuYEJTfIUrU5zLELaASQKX/hQG53f58x9/E5ZfjfsTjCE/AQSKxsEkFCi9lvBXi
6CAvfO2LF+CPDjmIr5wjbKpia9I9CYix06HGufCRmGbUmfdNHZDp/8TP9t1Egw6/MZyRMeXvU5Z8
rdCjEMVJGB/mRY4LPcQl31wNck1RDbtYO7rf1kOZHMXMmYMrXSrPltaACsSnvet3Kphx+KuoIfDw
jQINuSynAGCJo+0IjQ9q3GaSxlKfd6DJ00FqC1C3kZgJTAPdWu4cVLkgibhggSr3+Rt+yWlNyhuW
Ays8WSiHTm0S6Zt9ewClbazmpxOPwZE3LNoQQddpoSOAZPK+Xj2kEUwT2Lk7sKZwYwFYD0W865tu
wVoiy745Yw4d3uUingCjBA7WVbXHdXKAVwWiHuevAaqDM4Nbms8cbP7e2kvpmz6KGxjnprPt0BKc
F8AdEwCk65aRHodwzava0pBKYMBWG1H/xiW55MqkIbj6k/FAjdTYub+u7PTuZWCgD+t1UBgqlXfR
RNMIUfx924I3BWD8JYYbQ8uV+ODuDEHFSFBFwGdZa8ZKUvLarLQ8hSHVHdn37/JeLNVgbYytPpbf
aarPvvrx0zk7rcYccMFSYz4mlzQbMrEKFK0CGCmYrJ0q5i558GAPa7FWi3li5PgaXM/iuf7ndJLY
jZQrJjzSH5KN8QTr/cqx6az1U3bqgOQou6G0ubVe6dvbci98BTbHrW4txI0zORIGCo9tyTFz3bnk
/g/JKoLXpVGokK1rLQi4SRcSyMOo4py9LjAyKBeTHLBKbkJDn4EGJNzht1g+ohUuCnB72sxJ34Bm
CFUWpH7LMSH8iBbvRX2CzN5kqPhQNI8rIZM0jDSQiGIeEK0DLVng3Qd70ZVAaORO1ET2nZuDu8oy
NmWp84gPccQrruc1ZqQWZeBngI08wE0B3D8z3rBKfg4kF+XBeuZxDoH2mZ/1lF8xIY9BD39uk7ij
Z1EH2fbC31lam7D2M4iHJxsGggahKtSTxXog7Ikcm4TaGqnBpKbfnbsUgY4IpenxkUMSkF2obxY+
GA9NH02eeyN5MuBAgZL8Wot9cbCFw+2l7NcZHy53AcMmfILs9fI6CrJFP8tBnu6I/A3NLYtgDCaw
/K/zwtxTUmCinGnugTNKAHi9B4WyDQPnECKUq1McxG0BhsUkaXqtPOAAvtvg0sZ0fRGFTKZxzkkE
B82+gRK/Eri69aBVmFlnuyKEUYFI3NTNjgQ96WO1K/I7WhkN6TpP+Qa0dTErnj86utyFiVxZxuYX
ac6+0fAEA+iUNTpNFi+E2InrYZDUfwK/LMt2wzQyqcsV0OnZ8BePuMSkgsCa3fc+SnFwmpg9z819
9idGO+o2uL3FcX22W+ouURCPjxeD4qwsp2plBmV6xEqdISWPxqb7JHDT1LsZf2K1u02E4kYCCeKx
eQOUA1NbOZHcbquublwX7XP6kOeOTzkzZof1K50Kws/kCiUkY+s1QkeII9AtMs/CtX1T1e0h+Mm0
TpRXv5OGjCNt+011nMyWgw86gUGRpFYkMmiBCtNC8F+7fhzobwB61JewEOt0L2cUJx0AiBeYLp05
hkbn3UMxFBZP5KYTwpLmqJd0q0f18zCMmoks2LkLXjWey0OnuKiAGgqaW0B+iFSxngFGPssn3ClW
hmJpZH9gYmwyjauQ0LPjtejMxuTek0k1423Vppg/XdEofETMtjy3euY7EN5e7wSy3533Xm3RCKmO
jbg0SIxQyLGiHmYIKd4ry/oXfVgTk3sue9oNmCZyb21pNfg06ESPfy6Wnfu2oSrIMzG6XFBH3wAV
t0kkb4jc0VQbNseAG/c4CxfdUM+AAr9/zmUwgmLmYVXFXDoRtj2G+s3pGSY76LoQlubb1iKfrXfr
pwaNfF8PR4wiA/UgdEXr5kowjRMKDGw2a7It7+0/mbxW8ySwPsj9b1WfjG+HNU2VRsL0uFOLQlmM
c71lijGt+hPTVf5thpxT+Iy/qSJ9x7ChBWgG0dBoZ62mqHuBSnJ0qQRjWXsEwa0OrDfpO+6rmlqp
s9+yg+G2tH2CLyXh+P9ZlXKGKjZUS411J0GrKShsO5W++K0uuJHVrTaGKYW336vOKmg94LXLvmrk
/K7qnlV2gJU1QRMnKVUSMsxyvw0BZuMb2/2FyfeBHUW1pe1MKO8tTmdkXuwtI+X1a7iHfpSrJ3bt
U/Dkjt8mD4io+GuNZw1V2Gqv3GzkozlFvQZMkBjmE6m+sic+1WYWWigiB5nW+QfeHHlkqBpw1L0S
N0JVW7BmHoSwoUCQrAv2qARCGh9I2Znv8sEQ/RSsbd01wB1siN/qlItecT9ij4nwI79sJ71pN24y
P97igBONQagsKKfWYpkij9rjE8G5WeaJskcwh24fGmp6s6VaerPEoG5OiZ1x947uMUnIR14jcA4b
ovvi6JaQD7UoXN+6iIR4pBEqwbqY7q19oq7WVpCv21KPtL2UyE8GL9eMM/rNkeJ/Fvc1bnl7jlsf
b5Ay0IbGEmzl1b7JQhFpzbTROrtLDYqs8YDSwnDNv42acjGP6PgVVR5np1fq0JXwSeH4Li+GtGGX
A8ePiP3HQXCOOS3A0nYPaKJoRDs37NZuA/912BZcZzbQqV4hWoXH+FIMLZXZaV7E8fTRrd1+LCdZ
JG2yA3s7w9SfMv62cFwoA37NMqDs7ouevehgJ57oqDY/deEz0k9diw33QDXV4qjSZLKtvwSN7aGm
Qlqz0+B4WMKxUIReKxk6TjbwExywX3/EsuTvT0C6psbF9bkJz4KsB0HgmxgZFR7ievirJYTlxYFf
85QfdakeuEPW3VPtTY1n+15RWyiE8knTkGWoUbzx2CEQk9dhWfk+pEMph8TuKuuJf7DQJEan0qpT
8KIdHknHqhhXIIuuS/yReyX9J0Pfr1Y/PszzSFdOb/a/YWOGIrRxELHLPjdrLC2K66IWzArVO28U
3J5Jw5vxTX9oABagj35uJIWesLyTDFt9r2LKvjn0RLe7q0l9AUyF93Phfgjfxoeh/SzaX1U9wuKl
AHh70b4cgYplhlZoqsbVyt+FM9Hkle3yQU24+SzhA3HTCmG65QXa3UZAyb8gPaEzi/rsXbIvPysB
q27Jg6LOiDpMO2y/emN9iTW+GDOcknZVve+WW1btX0UExqlmWvr+ht7GM8zyN7zswON9uN3spyb7
rCHdRkRfTiPBxrk0d3gfe7VgbZfVd3TSfDRgKu1CMUp5t5BFYP2pzgq3FTtbpWP7R4U7ssmJptf4
A4NFKJaX9X7EB6rgXSBM3esT4GEccx0UK6Ol0pNKeyuyU6vHFzRLe52F2wtNuRXpU37WEiWc/+kD
LrbAsRMDhB1YMGYUIRa2sxcc9nNCOtiClckjEiS1UwCQDtxOFqfNccgLaNZ6OoQFyFpXl8bt+52T
ATiU3Lveb0x+exe5PttDOQ52UrykRJ+X8Jn+m7sFLX4aTvZff5S51rcJ0FBQ8fs6aJc6yPSaRj6T
DkEfeKersQBB69R42PVha3ZrCzjZXjp+CSWICWyGCIks8LhPbu/vXCYxgcY0dE0B11ucr8CvbPRc
KqXSMv8Tza4v1GGwjMnR6/NvcFP56ig8KqucGa/ZfEZs3WAyjd23/jdL01q9QS/YC9Yz7O4bdZFv
u5CrqQAxoGj8/Kw3fu2lZGzZyHjK6HRk/6IQgXL1bB92vYKsASoRioZaEx0nCAfYc1WNaUYWt2Zu
e1Gl9vVyL1BQ7u1DlBrUcY+NQgDJXlhOQMVRlercTLmOC/iVNhlbK3pntec2iT3UuMfXKX2RCMzt
+JjKVvpIq7D2dhmc/0dzYiNi10k+uwSPp61h2V2olR5pcu12IR7bF/4lsyE4BHe4jaF5Jg5skLAk
oeU5b3hZ1+/zcLn0vVUvsm6o8aR70AUsIlU1yBQjNsDWUT8mVMbpfgFtHBiQ15e8haZ3ypKdC45Q
3MmmKWlym/QGRK//lLfLGQAMIruqhDmvnlGIKI94j4bDt3a4NHti83A2XJiqBNWVsrotL2vSXgVf
GdhJvLZLgxa9rBNEAfSEQom3+fHL1YBZbcxDVXzq7Xy4wvzegcdGCuUB75iBeU9YC4WoQEkwjoXo
OOKBr0e4TykpOfIokLv8HiJWEdCxBPqNK6x6lPpPTqFdFiqiLf7HvjD1ATFRbtJ1tr/Ycv0datAw
/xWx3fnMmuR+y2yldQuUZzxVb1VXzsLhD6JDFzH8n40iiC7cjYcFaJ7x2opyOZN7wmQpigQE35pS
zh3cWOFgnGyE2FRYHAUjZQkCEsPJVPrG5DSzRlDfFznynAYEUJqW1CSPZEXRdWzVp26Q9KA5Y0jO
PhxRYVxNwWu96P8tl4JzwJUuyhm8GsQo7ObTTahEXIdpJU5Fa9Iu+mHq0lh9MEMkSqfuEMPVEkVo
eVAdIJiLHVcKAxbgnQFmcoZbeA9IsiTwi13KMLdMKYr7UFbBMaPcLJaH+BmL2+dfJeIDr7q+Fscw
KVKTOd5YEkAVMq97l5Z3evywOmWRM8uOPzKoWTKSj0FUft/uFcRiKq27EcJ2oKoANv0RzwMYaHMZ
w3ul+u8TmETTHAHK4jvhooou/BLWXz/HCVCPJ5T8wsdgW48qVG7wHhpmvwws5IbGpjWyZ0yPYZXo
JcE3CnxVfgEDw2Ao1A2Drfes7Yn2aO5DwrhaOOJp+u4kDdus7NAPpr0BODhKzJtrgPR1L7ThKpBj
JuyMUbO9leyBDp9EjqnzmXrkaaYqRdoCUW2CAyERj1cLxDVXGLcW2BB39NA3kcniwJ2520hl3xJJ
rJjVPrfZfeVCH6mOE442FXLpRdr12grq0IKq+UvTkFGypJONQ8FEbI3J0sQl0H2K/Ss9j2SBQiAo
TY+qaGayHvYPJoVWXZ53fZ1/mpM6RRVzrsCUCdtNpgfvdVlNlRaWJ5WPLkv77bCMG26mjEdHWyPl
/TJKLbXRvo2kftuTv+epQZSACw3XezQ+Os63NbIdF5D1ICFYqKJjblgUly7EBPKlLDYa4MKp1pDo
L5jSzwV8JK8d+AupfUq68aELVWiHNPTg+YrR6oR2ZUr+cPKXg+oGbTBlK/3gCwSKzafl8nnUrZye
jmZX09PMpYhcASZgXI1itFC7CzNT1DXFD/a0Semezburm6T+wesBTosgWhr/ooxWTNe4kBFCZrhi
SLw9Ea+gHWGwUu7Sx1xDr2Dm7ZONvO9ffvM4PsfNc5Lcp8TME1FT9LChuNiGxvyYyzxIp3auyYuv
f2z9clK3EYWmamjrXF1vtiMA80RA85szlqdCWj8BFzOTbakOLv82JdSJ0p0b8nwp9HjzpOloWagi
AiM78lxzVEdG8SkQFTCkQfR7YIPuFQz9h69jxRjvqi58PMAEWIm92WYEUv5Ug+TR/6xh5WWZ3k0r
kVOCaMHk8EQlp9rZ5bZvH/xl4JD53AIEpFa5Rh67nRCvBTrgll9A6IUB1yFuKspEnoOswLybHYcB
vLcC5K4Zf6DAsnhqyarGKf2cjwWU+YB6qNPpZF9Pxo80fq0Kr5o7/05xiU36gDSBhCZdXkRSN0d8
+iK748O2Jy5eAxglt4HFIEZg+nhFmIMyHhw/jPu5X8PK3LPciIEktiCSN4BeoFhCFowc7lJXlay3
ZsklcdH+++bBvZrGh3U7jguSeu0BaoGIPxPeWpjiEm/ClPNIs4LH7Bk7BZ2FMuyngeZyxV1TqNnx
NKx6E1dVAd0Bl8HmIzSGmJ0q25ys8H8V5oE/FR2/6dpXKVnIxpdXd2fydo6mH/I9C8iv3RzVYVSw
pbfImRUhRl1mxkj0J+vZzhlRUieivKiMolj9dLEGOm4WjB44zIRJr950SvixB3owHAnCcwakPaSj
xjH4i+aixXHv6kfx/GLqvosZD715WZtY7Z/BEbY6/t8G5LP10aeK+vF1/bCCLv3/hEyxz/xhDhdS
9iyMF3U1/AV/sdM0wtDuoOHqP2dD5nWblRh6oArAP3WcSj+PDVTk0kNCjTI7y16C6Uz5V/HrsrVg
XkV4PrMDToA4rztf7cR4qbAjWPAnUHAz8ReRZLl56Ab8DeiAOR6ccko8/B6v2JuRpu9hg9/d8T8+
LPqLoZ1f+kUqiVTkTFaIVFGbRFe+pxJbQrl5lSivHBD/71UR2DUnAybSg1vXqhpPVAFJSomLZrNb
9Wgj2cTvnCVBiQ5im6ppU+e1iJLkDFp26WA025tGisvVliHSIrnRigmT4lIQHhEDU7atJzQPqqJU
cPHAtJZGbiKeuzZncXKPtOULegTj5ZUL8bNk4/aecTCk5CXQEqGSlqtRSqoHn54i3QkzZvMTxGQB
mAR2c8ElZOn74MSrtGO+XoZk7AP1sRE1qeSnlY8lVs5z8MYGWUamRxWJo3l53w3BUsNBNu8A2PLF
vB66X+0rEsrO8TnUyOsUCZvZxx0F710R8WcPGUOM0y80nksm6GnYTGwzVa6mLWWiqnZgLmJn0sjT
vOLELzbWxvmtRBTqGno40NctfZJC9WJS8X7HxIDyJ2Wfv08PwsWpgoj6nofydJpvnnY/eC5VWh+1
Wxhdn7kxeIX9YUh+/Dq5thpmZSCzPm5yrA3ZMSaWuRZY9gyb+X8GBupXKISAE4wh+9NEQvO6KvFF
C2Nj9dyX9fHpzlBetw5bJ7M2gRBBWJqAnJo04rjJrkyD33bL0yjaigBLRDIiI0/kepqtMLxIL2dy
tH7QmJ33BEXxTs0P4ujnqJia3ytTT6fiJ3r/SLMD1vSaueQ5EJccXsvI0KmdNa0SBfQEJE/fp7tI
jHeXwZJXhLJwQUMT8PuNvr2ZNEC9Ek7RfttlsHLG3MDl2LNPO4TNr+RmQoX4dNWWjxcHN6+oQB5B
nvrEZI6/WcYA3jr3nAu+fiPqirC36jMHu0+27EGQMQoKoXjuRVR+cuA4vJKlhUo0zPaxecIFLolU
L3XGo3qifDrqIzoFFTBZ4QLhzklV1f8Sr8sB6fT4E5qTiApmSqW75GrFG5Wp8zufI8PhQqkMGovs
8mVWaPjWrsioAVYVeK4R9HNDM751AUvTNN5acg9VhSi8j+XjCiDBCx1im3lFkygLhzFzVT6BnNLg
X4D++wv8pvj3DpGwsPc9vMykWxiPmfsOh5pq4NiAfMk8vSgkaruxW94r91hbeNYswfKTmeN4G9Jf
PPAjCj+jGGS4G7jJnoviQSJeqhwGLa1IoZRFdo0NM2I+Mo+BHnve9EDF/hUsSAtJ1tefrT/YwpED
sPcVWTHeMQjCJOyDbtqknDf/kFRwC0BHz1ZZ0irgpQj0fowwehoPBmDZR1EKvLeeM30VoVs4ukeY
UAJeaXBThPvumE0V1Nb8DWYEzD0BfwG90pl/ZSaYMETGqKCYvc7JPY+OqLnqp7/4+lQwh0BCnsGr
t5VDZl5khR+MIT3Qwa2lURX58zwVT3+Zh4ufhreaJ3XQB8NgtEvohzEmhv5XpTI3HHGQonTLaPcI
qhUOyIQwDMfDyapg9XPaPzB0kFD73xb5gjEHi1No8Xp9rZOU4voLJ+5AlQ0KMJQZpkXpDjRgZQhw
jkXqHZDJT9puXDJG+z8ZeLkqjMRxpxM3dX161V+sInAQ5CG1PE8QvHg0LBvbzvBfirKrg/2GljY7
uSb9V+gbUMu50Bc+jt6D7p+0jtGpe5iavudXO5hbXXMM+iIU6p4jaMHfEMj4yNvBG4EBlyOODzh7
po0jswSkKw9oolptQZhbrN3TtDcSVIAPHD9XgrCF+vrn3cQaTGcJzxRtEcQt279MTxC8rM40DrbE
K7SFWyi13sFBaTTb7DIXa49FwDK2A+0Ylw6MFTPs9eILqmJsTg9FZDbeupVZiPEOTJJcZhZRTRTB
aB8GZ9P2pRz3SLZKu3nliTlaLaAAyzKjfO6FmKOcdoocyvOuWLqSV/QPEQqnz+UQPsnrazg/hBwi
z54tlp5gdjXTOBERdENn0e3Kp8ilBkKBnRSTuPswLw3R6wVDbDLvRohEvZc713veSO4RZvNtdUpc
aZjze0vYm/6k9CU3pD770lytJO2lMvIvfG1eemyt+BGRzextfyUUo4hOA8VrguoukvjbWiLekA9H
H1RbMjKm1W4E+YGukgv6D/YBUHVPetniPEuGJkbzKJ1lS6BorkD+IXLBFk7zxr3iqD4M4Sqeq4Zj
Av7Wn+0UOPT272Jvjl/9uuedXURp0SsSCCrFhcpGttPZsKCs97yuN7ch2JnYoV6S7hFBCkknhQUz
L5vS4aoMEvhWuUGqOnkZU0Vpt/+12a7EVHlK8blfBJHReVPXuT3K+WM5yr+WSSX7WUnyZkoCw+EO
B17obI2bVG8Py2ZDj0QkVEanwc97AItEvZX81EzlckssggdZjgeJwVSRZG+H1Pk31VCwIl15nOb8
HgWhZmZCFyCRHRxFRmoYHm+0Gcp4Oqrjv88cyY9PM9b2/G+JJHTNWYL7ftFxoJ9nnZ2cH3QN/33W
/0dBs3oBnkW4PA6EyBgExarucMVKbWA5PsOuLmLN+ncLmcsbme+1UTWxRLE7CYFTAZQS/hhsCWrd
RK5mgrKdijjcW03qTagct0mdLYdsaUsmxsWMAkZZ/dZpSXTL5REZgAT+iwifqakAd+SMKh4+gahu
5Y8GD13+MigaXyUM+0I8MBS2+uxl44TQCbcBCEsUiDU1aoznkA2z0ea5Oa/FdZ5EEjh3D5NyYzOL
UW6BMMuBa09RstRlrhuq/BRkv4JMNnBOjAxucJ6pgO2c97B7aLPmTVhcFMNLbQpJaZg3OVJOzP3p
YCJMZaNz6XocVpJszrkYLKgfvme+ZMYHu/WzaqJhu1DaKGsj5e7gOfcWnLjW3KE3AEgoNjPyxfqZ
tcgXoiSGmAZ0yNhxkt0XSTo2dIHTS63xo78GYeSntZnW+OM9tr9ckIkAhBAJ4czuFqp5FpwfX35C
mO52ETFpLKxzPM0ufv08xmPS/HFDurgTRLyaQYGHQlK7urQnCVaS9RohOEqUd2Fb1+YnV5ThkPYC
21MnF2iWhVmlgYGi4idCfZ4r9Jsa5lfYFxbJXVP2F87U7/xEyYQSKpTCXWCfiJjNhjR9jG0WVH0n
/Iy8114YnBfuT6oD+uMPimHITP+HPwBBIjRN96QLujVNNm6/LTts56e8SSt7QsoOF4Juksd5rPJr
n0oo2npphhWfi6VsvwchAZEbE3sxk5FLXHkYb0F/LQfVBc8SR/6UMTx78pMWVjtJoiV1iDByu4Kn
eRKqHP7dKvduF695z/z0DgWHIchno4qkD3SL1dCAe/X2wljaxt7xzDG4xdhvFF8+Zo1Z6fyMjLIK
urpTXsqeCMZpbYM/ZeZZtm2B+Y6aE/3mRzQPKlVpm6RoUquYBzwzkmoAh/zzx7qgpu3zYIyLQ7bV
UhT4Q4ovz5e5aatNN2Y5Ia1Btc7S4VcXb8Onc2QpAHpmFD3eXqin+jPlE+v3k5vREYUxjbu67rxl
mX9a5fLo7UhpPvNURqPRPO2qXj8pBYofmn4id822vhbrqlfBhn6l3wHbJDL8h2QKw2LuTWZys5ft
wvvgwwYDVFPFKLFPV5zTPhutPqXa1Thb98rDJ4R5RDmGGF7yvlrLNjfg1vgDHTgjZS/HfVosG6Jd
R0XzyEBqOJvEmWhYO8QtCz9aujiHsW8cCl7AE+Z0aa7202tEIIdKVB6U0VwxJ4UaCIQiIbRpWVR4
LRpzbuNO905lCeZz8TcDsSSRcAFyZII3Nn16WyRDfA1105U9EaI7Sv5tPbHZobYJOnU7WkbgpLRx
joLj4JfbkqSP7UQgX94JfMPgR7pmx2Cvb0TVM+avJORj/OlLRrngjJb2o7/q5h8HkHc6B2tfqGq1
0xZ+TPRfpv3aWpZxbQtqfaFFpSvQe+c/pnL87PUoEpRl2LRzeRz8512qc5BPPNVEpUa+BeIULTVf
Qepyel2/9WPmc7tawl4MaCXYCUdgq30yoqKaFHbYm6AwrmCvvQTdvurCo9otViy2+LolU6VW1pCt
7Qx0jz4pzeeSNvJt8vMcN0DEGm6fpkK8sW2ADcj0hx7VeHvFzQy6ogYN5wEusjL8gFgkMRrJb9Xg
hOgoR6TXusF2R0VQhXlekgTA/d+9B31HQFBS5lD/7RsijMZARglk0GcH0nAYtv64atwrGwAIzLmQ
gqpR9QNzWjJGd+31LL4Qq+4lGmSO5PkzjlpW9JKrkoXQBvfDfn3hzaPrK6Thsl20VkUQm/xA/a1F
/Yugt86zKn9hjn3wnRYJ98KKI/oPc2y7Du47CGGDpaQRtd8fyJ6yfHuUoQaLyhTkDeTjg6XrDAPv
jhUprfD/sjB6RwmWGp8YH1o90ojyB96Pn9O67mbMp1myPhX9cfO7ZiFcHsu4YvlJt9QUYnZ+1/dY
CncICUAtjSVPns2EXzJh39eVndM9heZiwf7b0y4DykyU67he1Fm+WqghhAcI07oflMkh8w86N677
rzIZDj4pSlkFXenJySKKcNPMHcpdtV6bkA9upjNVyx2jlZWb11jxV7CIG8b0sPR7HgmNGe+pcfAT
MRbIJckKAwBGzIaXS/ybA2jl9ZTVAsltDgOGJf7hAC5+9rC5elRCX9srP2yWHvpCsELL+f/Fg0Ww
tcd0Hqyf6hAJnngpqou/l4CjU0wk0DoFQAlLrIw4iwjuv/BQL1iYEskaLpRGSdFLrJIMS01PkPrj
MLLpcVWNDCjlo1nRUu+c3rhzYEPjpj+/yy7HiEhXLEKXJd8FvYvXMyqqaU6GEBMN1xBaQXdPOD88
rWFtUXoj22TclLjg5srSaSaj1jLd9/rq2tU/sL67zYZtYhKTArsB3fWAMzGMek3OmXh1ELNHd2ob
/RkghvhqkqwLWemc+yZ+K9/MPJGUj/WZyPewJaqeDZTAeeKUvL+xs6X8hxQp2Z+SvyNBlYY6Od6u
2XdcgcNHOSjZF5SHD7ci8Q0+gQbIHtmxOUlLhcWxy2BbJxy1InNCt2mBQAuRq3gzr1fzJSGQ/Xq8
oHU3YMTUW4gPsjqUOFClV9tH+1VRFH7ofCSyEI5GhsTMprSYSB0vgAgf07sihICvmTjV+bEpohzm
mYD8n6g5u+07B8LB0leHCzAM2AyWI6MoG98JHs4xsk3fkyDgJRiVEnK9tUcKO4Pf2DqsnIfygiI9
mFzzQPhDzw0G5bG6w5xbBX85HvYWMqwigRUKnzMe3Jrqs5ZWWCB3dcAPRjOk21mUIIOyg3W+eLsN
3KAHzEBNS4qOMDj3Nh3wAl6KrhSzChCwTdZgGqpJzOE7y5I8qQVpE+FYGqn1k5zv6bAESY5LhQoH
SHatlCYdRGNix+jxnVYk8Jfe4FTaZCOibD2voX67NHcKTA+FTfwEVEw1WlPQ/BeotVnnC9t7tUQ2
fwuVqtbHtCIecgfT5hjLD17UauSitEQa3oP8LYmzKImN8p3MtzIMPntDeHHzZLnDZpTso0Rc+72k
+oxUKyssV9DTNIp8aKvHJJjfGPkg0Fzg4ay555K0qS3Pu97yS8//5uSKpIgAQgl/NqBa3WjenffB
YckDP1SXuaTzgo1pUKQrgHxMkesu7vw1Po+AJJjqsnekntEIOty1skIK0NsCaXcIfmYYfgeJZVo1
BPtUP68nekkhm6/4orDieUfFt8pI081AaNdSw61x0zhp7MfK+JX+MNZr6j8/1KKb9UUCpMqmNOOi
Dl+Z9nlfAZaIbNLC0iI3xsW08rcmCFgJ0HsdmnbOCjqtVSVbwr0MUh/tYn6IngYefS9LmTg8/gaT
VdjjtQl0pN6qVhNyHllfJUdn4iS+k6fQlPWK7az6gcS0dg4q33qEWWE9hr47iqOh7z868Gov9MQB
6wqWAQ3GtjEJ65rYXhZHD9/WdT14bvdlAoKFyjYhO+L7C2aJ+1oNq2ifdifUwZ+DFyV2AjP9wNdv
5EGCZhfQEbaspwKncH0Nq4s6V5C92p21mW//PZHTf/h+EJoLmedxYu2h9l/uC1OGxhFWsd+t4s7p
sPKK+vjNUSfFRoC4+aj4Ofia3jBEI0hk/+BnbtIx6XrM5atpE0F7QUF4EDYhS8q+CJhDAHUQeqZx
eiFBbQsxNtDbLKQrsqhAGjlrQfViDG/WbE0CfLzIJ6+ASXMlc5MtWJhc7xvTaYA7vxF8Z1SJNPwl
aWHeqGsKpqsCGMW+JktzMu1R3l4fnGnYtfJ6FDuft+EM2rvn4NJnYnvTtKxlIZBkNTvup0t5GTpc
AXtAWABh72SlocEa9Vay8eo/dYY+lqYINQL95gnpNLREQJdVCc2vlIsh5Wj47we2ZRF7PLlhTfUW
FCOrQtNjiJ7QEk+V9HyQuPeIhTyW5Mx/+0q0aD+bxiQBITCqm7NXAmzZKb2j1CxIJLGuw4YasvUG
S6KgHdvAZO+Ddh8TzYMdOVv4rGiqKDYLpPsJsWvWs6Ns4oBetpvUTvZesokJplqJ5q3gzEBZoE+U
TkhYe/EUO4Xzgj1ZPPBq59yO3n1VMdKzO0qAHU+iuCVHoJz9HQX8RLujfy2M/kWodO6xEEl3cDZp
3epzz1anWePKwlL52Psu0Jch4tm4I+PG33jjD+sjHIgTNUfQE+LtLPWCMbdk2U+waGdCPx9wqv1Y
KbAwgiFnT72d8ylpuxjjz1Z5TfijCcqJJYSRhTivnUwIMRZyBm4osFxe/PLR3/eEGkDhzz+NCrsO
VvNO7hpHFYr83QRFeG1GYf0WG5t9ujoinL58KnHi+9caL6I5Ym6Z3n5Osdi3dZEJGV+OkU8jy8Be
nqah6MuHDnydn9kFrpKAx6MEAdjxZvaVz7cCDhXP124qRjJ3NDfQkDxN03uQoExvHGj9tiDsubCN
GKrcxQS6gOJP+6QOM8CWuayuQR3/khZtxNfvLAqXW1FwiRCCNoGv6kj8kDhhNe7Br7lmRDSMzta9
DFuY0Cqz0OgdNjTeFkZi/cffLjiW+5XCMJiDYQxsUXVH8nD3rE6jbRuH8Xhkdz6XGssx0Roppu28
fi8HnDykG2BhPYYMZwJK6DX1ZEN7KlQd+BXAZifbN+alPrCfcnrlGnjKYzALgIBI7Otzniw474mX
VZ0jyrO7Cc+ckDWptxM7/TOusEFKnFB6dlGtZzK5ReQJL04BB1erH9uyheKE6VoEnUr6irZLYC4f
lTb/4rlAi/Cn7JMl8hylNcPJhniy3nRIk5yL242GFct5+kBzdRxZCBiHnYC0jE66cl+da7Y0UT6B
YGCqA3Pd8ylKEfkd7goi4hR0zrzvU/tnrn+v03G+Zx2+MjauR367mQ+fXhsvPYi1Lr78vcOGO+X/
aOOSmtIenrhREHxxhKFe0+77BiKf/AaqSvaMOxU/rixaxJuLPMWQvFrd38L08VDJmTzngtHFXLbN
ay35KH8iHt4tNbyG23mrcY2s2xi6f9CMjrolkNthbkq2XpYkqNW1I4GsOJSqmuAsXkmTl0xhcF4R
7g1oKXKUfw/0+iaf8NFPBvxR3cm7tkkHRPBFtl9kcHpT3O77vtguQ5R0C7iQ9Qs+74DHLHvdHfPK
vzdXVzEd2WPUMqD+v6NQ6SUF2Gy8YBL1IgF2rK6LZ4lvlw7Si2w5uv0FhT2udxTPlEsLzwR483+L
w2O9kmtUdhtTIu9RZo/botS2UNPJTNOU2RTsbKGZA6+vAz//gSF0Ck4jGRtJ14zt6i6IRjWrF4jV
KnhfDDrLWD7tR2HMPLVzuM7rbDV6NJ+XeOojaoOYqmDOE6v5PrmVRb7roGH9fOWB/Rii2m3c5jOl
aiBcFcNaWmWcoOyN8i8FEXThkegmY2mxtAm6LoFk25QH5KEtq48qPeOYB+p7LfupIDTksrtFeBPo
2B08uX6rD17bvB6RzKLRwbIvk8lJniEk4uWYnvTSBtz9RN6/xCxdYp8SAv1At+jM7mY7TKTHvlDZ
ShL1DPwQAPNxFOmmTjU86ZyzC+m4KRLu1xmZnPDlF+MCHcniOAUcUslSSTjZd/MF2Mj4rBP9VRNP
TKOPb2hADQyl4yMglXr05/sfh4+P3vTgl0YudiJOTyblDXLZDH74oWM6jVekVqdBT1flDbJG+1tu
aVpxnQHjE4XsY5D3zwb+6j4XCiN2JSdVchAgMcgARUMwtyy2T7Xcwam/tnGjZuX8p/sLpJCqeuRr
fsg5ACy/REff9akGxWi/VYY6yr+YAJLO9iMGI+HBmI49XDQrzUtSV2YX3/LftiMYNYUd+OB6lmP6
Ky0gISyg/bOYCQljlqMho8E0ZUwXOHsDq+KapEiV83P5t3gxMJq5728cWhWclVLaOALbvGOJ56vm
8AtmJTOtrGDxLRzhRy970L2jczT1GweBkkBQleBf/BqdNFEkPNIRpYko0jc27AoQvRUyqCRicdSn
Qx4B8gPZtgnPb7/Bj8HhGxreWmWlGOubPjkLprs2JxR+cfvDLka6DAyaG7fF8vBLL+/F5H73GVHi
8pVYKHzHQwbbjQeOKhaxqI5Er3WK98uBAsEcewXRqy3PJ9lCgTfsd6Vf96FhkLjk/hoOCYHYCoPH
LE/cMNp+VggRvwLYJiKsnaKY2PJUf3zZTR7Tw2C6GSoYGwgjBd4hV4blRoqVgShiXcKdl7G1ZVgd
g4dPa5+1dAOr9dypww7Gx36DqgpIwHfARWlukKhZ8msb8lmNAvlIbrreleOZv/pAo4r88KYI3W9A
ixE8nf4SyA6nfw1u9nAB0NHgDf+xXHBc/Uz9TtgDIkrygoUqoydlth0+KDTFB6lVGcYvcjpYnE6M
kPXbG0AAqgPc0ZPSlRejYTitJGpaijBv605/vrlbm/pq1YumKNag/jyTjWlUAiatYrRz9tnexrZx
ds7oR+ij1ADoozDRz24Bmkk2LcNFUB7AzH5171IRHu8NNSfVX5KJZ5jT0imB999xhmuSIb1KEMr4
viczNFgcRP79G5NeWiKC/QZysoIoq++KFlFbacvZqF3H3oZNvRmFIY4x+gnujWdCE68Opg8wVAU3
X4COoLGaZzv2z+ZZLhHJMQALPgRn3FVIiIBnh7xlbgKSKY6HHCAhk5HXaZBrRSzSwCt3hb4XIJc6
egUJFmZ+VZyyDkzrfd+/iIwfwpyXnO1YIDsmL6J3AEfObRGE1UdrNwEVAMnxK2q956xVoMWXTzNs
x26X83Ho8IScmKk3L5x6XSJq7f5CPgcNfqN8nqfZbLVJUw9IGBKltniRqRTGYOqe86ZcngE7dGAf
MQEVsmvh64P63ji9VuXkTaXOWBua9EnsVFBX5lK8IgzvarfXlDaNG7AuOW27KfmmtlA91PdMb/Dc
1Klo9T3yOg462XBHDyHZuu8cLn6G4SzcI4XpuO8W8GM0k0DQlSDOJIhfpx0bl73JKjylxC5ZjHG1
D0T2OZj0/gETmzkSWkEyEeyweeQ9J5X/hyXe0PV5suTJBGguZoVKixcFQ7G0V9+GghAS6DFQ76Oz
BHJWxwfgOB46ruA4RxHuX9QFwICKkPhDZTMtCLUlQDqqvtTlo8ilGqJ02ah7TcoL5O6u/xVr4C9y
BQzCO6pT1viSQvce1XSXaxzS+FwzduVSFAKYhX2WrfdV6EhfIWOsuX7bJ7NuBjSjXIiGU8kIYoV9
34oZnyBcnttuCbNtoufjX9zoItpz31pGKX5AkZLgv1rdTXl2mYpehkuyqO0nT2+pLBcol9zebmCN
8JB3SJY373FN67phHQokK3s0WUwlEkKRrOJqEn4e7WufEOq6MTDe7TGGiAosGrhrmLI9DImyOHFE
ITr7kF54wRCborLCjCmvByUGdH2+5SVhe/d234ZEO2o2maJCwsIxufx1lLTIVe98KRZohhEwYc4v
iYRJeR/gfhdF2S3VtI5RjLq3uW1aBF+LYKj6jsjYfUh4GYYM84M1WFZZAP7yUN7af6t4+2Jm2p38
UIOK8nm6WKeGAbvH06MbeRGfk/xNFuzZcAgmUJ+QYUlM/ydy3Gp2DCnfH2XpUNt693kVVJop4QR8
cGy66xZfUKuT1qvMF+DxKzS8f7nuPCqx/9AnTQ1ZssLfwtuUQxybwUmi9evOZpUNwktstT/HndKT
Kf1GbfS/Vazw835AmB3QwDYdOD4jowLHFb7xUNnJxfgThr57WeAMwsDwR07ftQRj9TYGymGEEajy
cMhAMcLZocaTMERLxurl+6Nra7J4Hs8XSxrwEFQsPMfjvtEGHe4296RK3Z5jUaeguGoKPzGWyG3g
ggV0KKUrhNQESny4j2b2Z1Ork0azZY4Ea/9lmB7N/0LCm5orKCnoW0LadorIIAPoc0uBqN0buyDO
tI2703b8A10X2RIlHZz38EHegnIKGppUKBvbUGkI1a97Pr5pRrdYLcLjLRHHcFcTRDNKIvvmZ5Fe
yGLC83bjr/cI85SnDbPDutWFHuKnxDyJfH0lnYRGXj0FJjAx09sB4wuclt+IrwCl2yXyI/EMjs4d
P1T+BBGMZuVe9oHhd/BNCX45IeXXVy03mi1B1ht+tt7JB5QvcQa1r7IPvF7VytBuJZBFUHqgb+d3
zbRcyGVA8KUzBOVZdw/ReyeGza9d6i+PzHbFoeWWL5+VW8SKm84IQpx2NBn9pTn8/MXh9uZj7lEB
mZFskFoBZOnwgM2NjwWNjkxwoN91JOSd3eSF0nfJl+eLiT1ur9Xek4Plp7fkoPGMiyDKbJIGxCRb
U8u7oQ5eaGwxdeXWvGUI68G/BRufOcCU7SvA+zmPawQMQs7LUBXeqmesJ/Nsb2+ffBbRRj7AQa+X
Vf9aBmwRe32CABwSfzLWH+vUmkwxPdlM7mX4b0MpQDN6EZDEZrAsdliIG5rx3hNt09Rn7l9b3X1N
Pu8c2NvzsXAJAePTydd0S6RBE2nb+hoCkz/AXd/q4b56e3iEAAOPk5m/6/YgX7lliS+2wKF0P8Y8
r5/1+IE4AFqrz6HBazmTS11NH5LurMejtCKrHXBAoB3jiJDlk7O5tOu3MiuN3QRCWp8rcSdzQ7m+
UEShBxVv2SgrONSSaHhefh9zJE33ICf+oJIkHtRAROYOmr5IOUoB9US/LY256adANc5dZef861vS
wMTadyNR+6VxpPTS7p/blV9du7AWhNLxtGFY6obr3L0W33MjQthnqExsUfjF1eAwVMrvUjw+HGQr
pugmkI0LEH1Md5yiFQpCv171dsv7QXNvNzItlbr4KORGB2WGsD8/l2PlyNGbHZZJLLNWQygzLR8Y
yuDdCqmWEOaMbubWE7QjzPYh4idnGu4aP9Igv68B0/AS9UG56qmYIA4lSirDEPhzO5m1emNmYZfA
z0D6snGJimRB/Gv6L1Z/AvggaDs+WYF2hmhosAyclMlTioXClY17gz4GLoJ9evxIBTHWVlboI9S8
fidaOl74doaurt7+ccBLZQ8lH+RQXzK99EbABO4kvYR+azxZqPF+66Blu+rAyFTz7OujPdkwBFYE
nQAYL05SxWl57AfT+Wrt/T26B+fk6ApaLU5kw5lWWXsiMe++aVJaNKWZFuxag/1dnDWpnso5dWgI
xDqR10xzJDd/Hc0wriz3M7BiXfWsPDgzyIZcLkyntUZoiJg5Tu5VW/8tWX5cqkpLVt/sSV4V5o90
EwRC5PDTXcz6j+o3wDhxvROboeXSwErhp1SEKPRZ4Er1u4HiJ7sIp7ySlSePXrfGS5AxmrSCUW6g
7qUjCs9WVTjWhYxK3+ajuleYNJ5CMRo8cdnRO4p3qigeol3ebCS08oSDOjvY5jmHInwPI1QJkQOB
GsoOEvTWQUTQMwA9bRia+A7mQkeIRa1s8BSSWHqshJzCk7CkZdQzOw27DT4PWtFDE2R6dXNelfal
uASrtWmd5mJ/Mc8DuM0QAea5EQd/eLrKafvdTnmqEHwK8nkFZIyaYFkxD6i5PMEu1Wxk+sv3byh7
F0yx6mkjOrkJfIrffczE8/zgO/vqUcneOj5tn9GQe8TMqQicyKhr8hDKsa7BqWgDwf1uKMLEya9Y
BKuQTroEEFPmL2H0KYDPkgyKVk/BjZf5iHXhZROFsh7hRrDYWdNecEBf8hx3mLqG9MO4OVzc8CFc
KpKOKEAi2mRGxLS7SLqkMJqUawrCfx8PooLx9T2w3xM4j9UNOBj6V693vonIVgYB6Th+IEhbXEqK
Xh1fTxiuCdFbB7+UaSL0zGm4z6J5W5/KPYjP6QrKaseOUHkV7k9syjSa1ftAJGpmawAX+e65RcuG
J+57ZHYJa/v50AD60xV0xvsvoPjK6W/Tbw4prGgXWDJ3h+L6kAMfiF2+fiLCQw+BnyFV23Sc9J6Y
fCLkAq/csVvOM419yd2VRJU/IlYJoAMinpO3EwIhuHFyLNUR5HrmKuUmmQBFG/5cvIPbqT4SqY3D
rUiTAfTMGcTAIqi7/QPNFIz+M3P6+yjVBoROB/UzseNw6eJFghvKM1WJmmkE8E55G4cXrJyzDCjX
TlatWSvLvM8KhXzTKQao52Zcq0qoAyO20YR1Jl9jkv7KiF932Rurf5VMsM4w+sI2Wa8KeerwnLjQ
FUItfMjYp9NCYV6/6CstRA1xZTsykFEcXHSGN2SQ+Xqkw0UpkG2lMd92SBsuld/m7Hzzghm6OLwd
RXuePeYfZAiMRg93BlyS38ddlBdR9hDz8XWy/yOBqgbrjB6ePA/0VQ9nverd2iDfPk3jhwBbt3pM
Kql+4VBN8mA4mxGcgX+go2ZCFKrpP4Atp+YksAVzFJKaaFgcFeNAnvoisPtZpdttiSYgf3PUX3O4
l8BT+NCalklfgfXaDqrPRyZqZvL1l9Pyw2SzcROUP5Qy+Ws/W9QGTpRfT9IPd6EhlNqFv4cJrMwz
W+LuzXulGCPJN4AcmUYbgO95DCHze6jBfSiQYpFJI1pEZ5awxpXAWADfT9G1IGU4WU/vWyeDaHKV
Hfa3G0og03Nk7MTXh+RCXXK7agWdb1tEWKs7x5DtnQf1iEcjGVyiTjxdOJL+KshiubOSmkRu4pGx
mXGLZnpIOFat+cyl4PaGqPU+ijp55HQUzNaMynh8c6jvGybRrByNCGj1HEVwp/n4GORpG1UYkzRC
1XJdNLmGjOzo7qNYs7rmak4RFW1ALVVoCx+22Ca9X5X7uNAk3O62l6EHWToxIE25IcRJQEPerNDh
WMc7wF89AfuGBDvz8jjxjEggzG/hhaCtf2dAhYDt7yA1xa+pK6xZwYWzODy5FxAOSkMmzP5B8pnj
GMBMrGQAZz+Upx494QDbd57GMAUnZrGcNvhSFbBFJm+LdaZNCbeWFWQk31clt780qpYQ1Q7Y4qmO
O6oeymtzCn+u4LbywXONXZcGRICpeUrisEJTjN6gsSuEImNanwRPGuW5o6z1YifYFqqaFe+EewaS
15mWSscYAa0cR1Mw0BkVqscigk6q5EBJVh8g85MdB4+uqFXKNcsLSmUtr6KlRssJAMTkGzVnjDT/
du1SAlErnWx76sNvWTgF3uq+IV4jc9Z2D/mO3LRGckWqgzNCu9bxXHcWs5OV+88ab2lEJkPyF7vy
Gj0tqXWqcPvBSFffPh1PDjDuydNV6Isb3gSgI0PdX2M1KS5i3uGK39wWptBpj1cN+i9T4iFunNDT
LybdhZ90rfz6+Cmak296XxYy4hm7StsoJMtjMap0ybhRDLjZ0kuUG/oKXmB/43R2GgPsW3mFRHZs
utZp4wFuS99rreEpnJT3I74x/l1NLMbjU6knnV1797aw/++vTzv56sm1RkjZuzHx3EbLhaRG+WUd
CfFgjlf7mdZHGtFARxV70NbVs4Ta9oT7iwAMAzJL57soA1J0zS0siHM8wwazJGw4sdSXAfTjP4eP
wjrP7YMEogqO0oMxMSjP/PaEbNx1IBQlce7dvF9BRQdoNjXipPedljN7/LBHL2QphKvTg6MLT71/
AG1p/ywai/eVaJHEqk1GUTDOenbF8yL5zSlV0SqPVeSkT3uPWEaC7YCHrYJf1RIaP/SQ3ON+gJ3F
vOnJV4VkJov/4O1VU+kpOe4PCwiqpYgivfwH3fyB5YcE+eOexbdsw4jPWQOlPIlQolJ/Bks9/jQJ
dyVPshhyx7Ow/leVETblg1kJR/nZLTCpuCj1B5je6bQsdlg8+UnvlBizpVs/0+ms9AcX17rqotmI
6HhC7LTQo/T210uORBzhEs+gjdIDS/D6iXKbkhmg87RvYu7Ms8TF1+IxjnLhjzMG5V4zuxQfJTsm
Kr86ngSpjs/iYlE4wPDMmZw6q3REHH46kE38VueO+sLHSiS6sxCs2INehTbBU/puCe8sF+ZUffB6
QENZAG7Jf925jhr5cKvGo2TGBR4jNaX46f8trUZqrVevaSDhgkiMlFKPllelK3vy9Kde87cU74MI
ro+ltWKvR8rWhsW0/meAMXSgb+d+qeL4qo9DNtuZPkWvyS8FkLl95azkh4clqePpBaI+2YR3utu2
ncaUeJGnjAXjiw7eDJ9E6LhVS51GVxvzAZWWQireXH1oR1LOpaqi3Ux6Rl+bl4IyrG+yT7MLeePI
zxgEAaCbD3x5xcus/HPRsOtEkc3pRSj8vO9s3V90CqR7joHXoVfbkE0VfJ/nhq2b+ymGa9YNt4AA
Cos5iZ8vzEWM03jDmilVnChGh8CiGePAIeAVD4pMeRIH9hU8E4UhO1X0j9gbNJNAt9xUmRMgkPJT
JNJIQouDRoq2/RAkEumqLYC4lazWsykBxrejVIxe/9ruPWbSrThMpp24wk6AZYb7okymAnTrsG7a
5EJW0fW4AtvH1bDi5ymTzqJfwonxwq3ReF1dtJ+rMahihs1HyCdkXCHJn0z76rXtBEw1Q5B914Pw
qGbCXbIMKPZMwbyspIQxPy1i7gt6L6kyz+umCiOSwZn6CNy2GTkV5AvaACpbuD728Cme9jGtMtTP
U0MpLzClEOEK6cOMWvWW46TrKW0stYNKtsXAb2Hd29/bVbarbmBkmrjoK636qw6pgJZLUXRPaGrE
B3CG0irNrMDrxq449i/OayD87QzROJDReV9BFdKJfWwoVgkwVIpT0A/aMWdBsjejLVroBr5w13sP
Xo7HXhH7SUB1vsFHExuIUgNLlBFqkjkqQuVFxEOXEyaq6NJdPDX2Ga+83np1dPDnPUwJ9m7Ev6FM
6FRCLAZdC+M9D6O3a8LuQq5S9By+Al51SGz628fyu9sNjK7nxjwdR+jsKAgJqzW99qWkzeK0sAE1
3R9ugr+i4ZTDaLbtmOT6KkOz5DIyB21drhWiKXjiK/qNnfi3gqBemzRAhVgbp3/OEtqFoj/5Qgc5
Bwr/hYbweSobKI2lC3UDYr1d6N7A2PvHR+REF2OwErt+KgcddoTc1ChcY9QrXz1v686r1eol3AXh
N7f1SDaN+D0oKRNm/eCENHwFH9IOTfiWP2ek81zxi6im24OZI2ZDDwhaazSYbPNP2W5wXSKgro56
/b+FfLKUG9ByD6hE+WS1ADeC+jLQY1LGXmidb9eb1nylsjOEkRGMFbRtF68JgMjSWQSLP8bzqpEJ
q9zIYun8k28dhMUuHdzotXdNYO5JNJ1dnWrDqf/n2FHQ1GzDfcRc4PQVkcryp8DcR2S8dTmi4NRk
qzHV2PJCXEguFWkF7/Rzjv8pO1iwaszuNdihCHwgYIilrdSsBTgTcpyMghjJpYYLDIg78Vlh3zTY
5lfdhNrjlJtxntJHPy1gp0QzUiUhM/WWcjHhkviTDvvVfiOJuc/EAuIvN/IAGARULBcWWmR0LorJ
xDu7B8I2R0we3gU0+b7hb8xZTKP4DXIqu65KJm0lDqWcSRuOw4px4j3va8fiyr2vIoqSqv3o6+ZJ
s/4HJwH/jLN8iRWTDqXcGe6eiSiiakRhDadZLxC4m+Vm1On1uGoMq7rdpRWU+/qJIBd23TJloRlv
KPHIwUIOK9mOjabW3kpu/YttleTzEzTQefjcMX8uSCVxIfFRhy9EJvZOG4mVHu+BqVjeaQG4kbnj
K9upiyHjGOU+tZOVZDGwTR8XIvMjSUEGQ8BjPQ2vNiu56E/zjsr/kG5AnPa1/fn/apbuppv8N6u6
4ySubSpiJJM8MpDoJq3S3ANh2TwjVJu+uLiIgeX1IpvLuTG5I86HR0Tgsb69smm3qTE2cETajaOf
1J+EhvY1ajFFKQuKNy1ncR5QagSTsyhGFrPs3Ih9rdtv2mNZPhnK0nPWtGgEHkIvIsDRXdU/BsiH
esxt9QtT7YPNMxOclul/rzhQaeIoiSq9a0Ub/17xpuUv3iqeSAh/+JLGkqk5vTf70BYl6sBXVmUS
OVX1J6IuMSC/oF+U61X5Gbj6uCH5chefc4hazweCVoNh6RE3xD720wFPSs0wTpfJQ1EZR/GmPUAA
WiWNK/4s8FEU/lvVJ3e60tP0D2uByPmQXwB1ZMd5hQ2qAn4wWiVgP2ngtU+Q0KQVVUsvMfo6j2c2
fhtJGWrsnLXVs4mLtyvHFmVdpVKDHvpZNVTR92k9g91eQ+CJ65OuiM1nPT96WCpYWhs+OZmEN+TG
srTIElAq7cFNRR8dhsqK33yZYi30AWqBpcQyiYHayPBhguTWcynptLJa/AkepJSm8Tzwe4L7XVWf
EOmbbHOCeKVJTww8f1R3hyGSXwL7vmylpl5dvHUnT496L9JdEyxMtzFRRQ3fjuyEgHI28qk5tNgs
ERxTawuBSjvBG+Ex3CSdfQ55lafF1Zmghvuy3VZVYEDjonWN3c9nX62L5Q96rlJfmNKD2gHEtQaF
Z/JWLpWiklNH2tv5FzUadkzQQwHdSm8P/Q4tP1x7Mpb9JOPoejTyjVlBS32rxzws3pEq8Jzp5c+0
P+uNf7Msyx9MwaA2Kuq4QUiWk/6qMaxo8gJTWhwM7FqBJdoFC/IkPR8v3vYibwJOYgBgMRApCkAX
tC2t6UGVNcRcWwfMVk91FJKxXnpguffOMlQPHAOolq1B0XtTs7OhB4TT/7P/kKMTDIZUyZ2me4nG
b0Sv/x8V7I5Rp2h1VtwuMm1wq6z9wKVvqzDey3LcmJfc9dG3yGGbenTsIRyIZZ13MROrkrjYquPQ
obVGYxNjmG3NHqBU14RYgmGa44QH1NPtSMcbcz/pF7lOmev71jAPHEeD1jXRcWFYzS2YeS6yutYb
3F8FyvBmWGAQzgPYG1DxJPNL7pummY94bRIfn+NmBJ339tcKuyVn/WMUrIpP6FW9c9tdXy5QLH09
aTM7GHFge5Rg4ubuBjvsd/RTy7E0ASlQZiW8OR3loVf9WTiwCmNYWqEjUC9uYUrNw2zvuemMLGr0
YQ6g/isZuDmqv8NIw7yUBTTnEr+vLt/N2jzfUbHdv+MaCmMEvNXT/kEaCX5rQJOEx6nnKXxQRCfn
Se6IHZhNLUch7DLIW5lBdUawogTrhnqPQHtxbArEuxW8ZfbIV+J64lpCer75/a10rfRnScGmcHGb
2wlm+z0avuF6NbEH471blY1eCqNQWp17ni+gR3v2Xnn3JHkJbaUGLdcovgUCmTaeNJU1V2LXcTS9
lNf0rBOvIcHu2JIErOiXgy99pw/pc+atksAhLfwaCfOJnjt89l6apba0rxDYMbyHUhZNVi7Wmc9i
VuiBs92vYt7L/nfNQBjqCBOo8jhhjUM2ZgwqXpmMf1OTjedVgyjRSS5dsE/g0pzDJvgfMojsSAkO
aCRm/jNG/eei53SQl00xmpSerbgWdS0HsOuoIRZV3d86qLUabpjHgFGWdMbw9oMlaJgrSERreOVL
siQ3nWmYoTrPnlO8Jb96ZlVgc7xXfuZr8ypZIpjvBUeDhoihj50S4jFMBln0XvDNb4+tyhGjNpez
r37yoNlywi/Suxi5ws5TJvjX9mSrm4QjNDb3LA+Cz6H60xLCftrnRAeg1eQjndLi2d4vFbmScU7G
cIbzmm3NOrlpACcpGbfzpPZNM0MbZrdQmpuxpgcpt4e0NGy3a7+mkKLuRoY2775jE484sgqJyY8Y
Basld5wLXghzpm4cEWWlMy/CFFWFNJGg8vHfpU6ARRARhgXQePNlFN3bwEsTkq0ZXPvC4OvIG8uQ
hW9rGZpXnZa+Ut6Oqlpe2Z8W5cu6WXN15PmCg0fX1m99lQ6YpCuFFVGrBtbTzGt4uaHFNvSr6gKf
Eh/weLxQyITQ1/Z9VYvAZRq9QGRZWr3uV/X76fPFPtOVKbKPiDhNgT1JCvOvAVL8bkLSM8EUPIfN
eIbD8KifMDgHy5oVy20j/6Lq/+UBuu8zrQUz8eH1FwicylsJbNp9kEeEUR9UuCUWD00Ka0QnoxKs
lqMLkiNV/gRgjfUuYhzKmjfg1zHdKb5D/+LgSCDap+Alq8MbUYl/fINDlFyYMelZmgyv4cqqXhuR
s3GNNGc3iT3Ej8LSoXdQZeYBTWJlVXb1bcNusRpes0weezTrlbWzoL8A9huI1Lo/Kmi/FKn2lLEw
OBh0YmpoBfIQ5oibQ+iBZxbf5T/uN9VzFuU74IpKr/wLF6uKFvdxO785fYozbhT5/5R89BZLnhH/
4UIvuz3/6SP49BHwxUQknQ0+cEZXeX5bJhmrHAW7kzNLab47i00QwAWxST95IhRSGW1GgkX5FocG
9DMZ4Y5XheJg82KqtyovjbsLbpQq196xNSlgvzwhYWhNBU8F+KkEhVRutlh5l4mWKruX8hHZ2C05
mYE/CX9Ax0Uo7QEZey7BmmubsxjioPxDTI/7LFH/yKTBmDxXeny4QESbGwmn92NeuadNNaq7aO3/
7FcVDoDsrpETvMkKc3o9TMeq5vSpqcYtELYZDumjXwY/ZgNVknfUf1hlXQtGUriegfKbYB6pVDhZ
YhW1J+jr2JU7/CPDOaAsiVHyZgHfgXa8hP0tJEL1TKO/Q4b0uou7EKbzWs2IqWEhgeAgEUpzTw3O
e4PTUgarihi/GfmPzH4YTG0B/nnnYs1yWvHim614KNWIiw+LS0b1SJiUMrKgx+VvFHJpXF7MO9d0
lQc6E2vrMMFtkWVGyZUiWtxITGyp9pXcAqTs5oOrEZslPNFGOIIcY6grorZvs3QHZ043RirdS23f
/dcsY7sVdWORUXMP5Aizf8NbdxiAGbJHjt7g8vzOzBAgR2M0poXbsd9XlpVlo6NltrrVR56iYNM3
gulxc5LeKtMuopgVsfslA6W7JJgFAz9LrFp1rvSVFQrATg+PN97j2iMBR8m9/Uys0roIaTXu+ryx
yfOtCEPT3KF2JXRTXH2rEhCA5pEnwJhZOVoK2ZLiyE0179wl+QJXI6lWX//Xuc9i0anXVj3yeRsa
dc16KUjh0rAafnyaU7tE1bTzQ/tFbE1YJxIxDYYDF4vUiPo0vKBzpzNizFuIWzBGjggPqxG0LE5k
8Df4Wv51RS65qIk9JMMo6beDoVvWUfzcIUMqQEriGq+fNiF/9q31P1ZVcvSSlfdj1Wve2ReHXyRV
DGH4WukY1r7+z9D3PcWo6vDct9WGT02ZPne3eriE9+P+vdFsVLYvf4Qft5HF6ouv12l9vQMaAcqG
hMqoue8vcQK4pSj84gu9O9k5myDM0K+3U1wXyQzgNHAPMzzqoqR4rQkWG3HGQaHAsNXRfVK8shyw
Q5LVC3cGMcnbfBxeBWwSt5q0lwwk/MAncwSOe0lB2V1OrHdy5zgifY0DU98lVKkq6vqYU4+DaRBY
q4SMEscomxgr9arkr8ilfsJ2wq7Viy3oRGNxOSIRGy9NvXz3XJoEWzjD+ys2QrGHHkB3WApE9M+2
+GMjKx4perKwNSbU9CI4vwnuI8Voqj6v6JBHdb7DTUT6rKfbKbYmwSf8i05SAdgEVjrqzsxCXse9
ipf7jlFy41VNzEYWB6+MtlDoS0TYtHfUcWuqOsnQfBu9SA6F7kmHISyvRcZkluLLKyWFegfvaamF
3PNWb7Nc9H3m7UQVGLDJ9i3Ji/bBAy9zxTsze8wHJ2hgw5NBtOZNk1Jx8kchLnPVm8zctv8TUbyD
bg+diLRBKwQmVRU8ZOybN55XG4VJAVUXbWEPor1V1GVyZCrBUTx/xVld5karTzdfB2j4VCjF3yMy
ECG7TZ9JTDcuvnSq//9ndFJ9QNEpBn1kDdPsTORVymQAQJuEqSbz6YZ+4FOo8kUtTAl8uox5Z3Yj
ADj8nTMm7zzCIkSS605EpDIChuXk6XxtBdTgsIz242H8w3wju0oN3qHQBStENV7N235+NeAoTk02
pq7smTZ0Kc6tfi2+5yz574WM91cLc7bfhjC1pOdeb2q1x/++sHanPvILlX1sXLaxojLUmBsKBwak
dH2HD5ob1UtQbMfWN/1FRkim83B0FcQwmR7H11gEsOFzKl9cGfirqgiY/yyfbcpDN9lpen97lED0
wrmtv1LaPbEptKYhR4nw6AdC8Ck45W9GGZJNjI6cORgOorT8ZBltEGYq22Re9o1FcXWfowBe6m3L
gahYgrLPqx3Lf8gZ7Ur8eq/YpTzN+n6cRMRjJOAGPI8H2M5PCxCKIHIo6m0MHh2ozMoka3l1nXpH
cb6zyJ3V2M9RoX0hpB5lI0ewzw6e3u1pD73gxpSBEwApEmwQyIiHHm5CjFlE8LPw1QGxjH2SQNfQ
z32h1tRFMxQBKCIgpKIxJf4OvLJkZwFe/VBcWpCg/Otv1jn7Wfaughguqj5cmEQ8rw4l4aPNAhQM
D+/Vgfbl/w9RvFuaySnTZ5+NHgET7UtsFcHJUWQPMNMjhxm2XDmiDhDFOFCrk8O2AWaOzaQsb6V4
OS2hCAOblK1IZeZCUe6+Ntf/gyMlGMXavH45U+xXW2Ii+ENX0J7oUs8rHC4gF9DgML3M/piuhbUk
QDZrWH9QWLo0aW9xAIFEloFFjMwAIRpFePxoecur5I/hDn8vXuApPoiRAckCQ8zSwzRPq4CH9+Eh
OhjYoA3O9PS6cIhw2wu+va0rURavNgItx+thVOp/mlgykWjjSGPEH+uIa081gUZxUiI0hJnwJoo3
ISokSN9nW/6okpZv311ar0mq5NfcjA6921dm4acr0AuFcDWYdXPFcOqgRN5Gb8rKJkVcHumSM/qp
n1Hrf87IEkhW9AMVtRDX/816TC7WXdpNfsCvBbvyjRovQV9YvAQh0+Zg7dHdVbY+euknQBT7wq8d
XgIbWtDxWl3yI8bX+qZXgFEa5rIUfh3zaU0KVjxZrRAz4PYat0Cvh6Yhp1lA/atobibMhA1ywkcO
zkF+XV221YjMxgdiC3dijv65j0/EpsZb63DQpcIKALgO6oEYhhtidBzHJKYtmJegwYiyKll4UKsR
ozSsDidXm8hv+9p4gnh9jCANPx4C6RYznyuBuKOw5eVzmkOMPSEEzXYfJr6q5QLNPd73on+Xeegz
PsfTjBqBQDrYWUIWGmCeFX03VNQhxU/lyE3Tqbtrt5O3Yc3NgRujZGdpQkmWuEhgmunk81WG6YFH
1jySuKRnLZCi6nq46hUKXjcRDdZnrQP5x+b40ja76FOh2juJ+GTlDS6CTny+0gT0s6o6jiS54ve0
+3Ilb3wNr8lROBlOsOGPB0TSl3putw8mOrU5MAxWdISrOW0cYNVUOkqY9rlAUVyIS2tQk83JyJMZ
hDKdI2hb2B83LfCmdNn+NYtePDVLqvFWALrH6cIUd53Nr9sj94ZIVy1JhMEx+kR6iQVDuSJqpu02
D57Ut9g24lhdrcumuYjM+cgoGcsT47RHrpgsa7ttlyeZfm8+qV2Sr0nKCcHIeEFu4OjtvYsyi2pI
5bCEFRPVotgRlYVjRoPfq5J0GJdcrghXMYJVDZMnPlv0uhUReGWQuP8Xs6qkR+XgJs70o0AM8mWH
VqwxLJuh9NN9qpIz1zYH/LR2N8sOlKDAfYJpWb/Ht8sGZ5Zw7FNz15+cKpPmXCp6tZ2rgDa/qtCq
jSay+qOmzARe+ZT005JnvRDTwovT51bOxZxTFdrIYh19hzgkU16AMtTClLnxPdDTE3YswS3IBJDH
x2/FoAvXWm7hJwUWgpqw/f6haKzo3WdTa8uU/es5EcjXHBCxq3ZNqUqUORnf+aphcVPsk/q/vAOB
69KZJSM9LJTVPb0n5oQEs1SabgrnOd80mYPrFybvXE6pCjO/SBq2GVAe09hlJT8mvuEJgY4mKuqI
Q4Qq7jixVcGATiXp3hgzSXk29sw744Fc+LYX0HCaIOUUIF81aQ//P2fldWK8LmS8dX+UEcQmwhLD
rxrM6Ic3M1neN3egnNoIrjIPlr1qDVXpFYKkII9we0h36kFJu+OXR6kUDauoNPtFiDN5P5PwKAFH
m2jnPAzST+9yRF6JTCKiRFPWWae7NjGsoZEcewuUtuhmsRf1pMv+QU9joKQTsx0sAMj46rmFG83/
DXWginLa+q2Tre3baiCX09R6JxZarqNNEG85zHDjjdeyK9OjVBpBwolYtzKjUezX0TaCNdeEgJ/m
RHUqSbQBq97uN0xn+zl8Q8cB3j10uHSOTiUsXWiY2jzELUC+yBPfpGWJsq1XiUfET5uAEK4ci68S
F3jnVtEcw4fsTfQKqkocpho0rXl1mGNalo7XrJc+g1kF7iT6gwTvOah8C/PGOqUTXdhxe/Be1fMC
3Tyu5awpLuFHS/nzzA4YhUx2VZp3bHNiYCq1shDjNuAdVLpVJJzm0ZPlSQk07PGQ93om3XsA+xuc
SbAft3q2Sv0FWIn9qqHYeSM+WfzQbzOSx0EtqTplMfQCw74OyILL7znEQ013FpBbpP7M01PEaRwb
5K00qmpX1G9aAcO2RAJafnDJYHWpR/S8GnHN2Q7a+0sa4bWLQaFK84pKrYkVdz89TKXt8k4+DZEz
zHK80ohwnlnyjvCiiqaofhz9hADS/PdiLkVRIKdvbbNm87/PKaM0Q9x7BWCoQb3aQk0fNwroV4YS
CEl5t6TOT34ZxVzk0pnvxdFUn36QhJ9zs60poYlWIguD7A5W9Ke4YRj4BcUgGhs01zKkSavWnBpL
TUsSoX4aD2+KU2F65LXu7WKOGcQ4j0nV44r0tmgN8K+PsUAJq81T8ehI1vcWnyt3Rb/Pws1H5EJp
+IJjOajGluLZFR5tdScs9dLZNnoAHpKRIsHaiRfNp5CjfGcMbdFZLNk/MhhgzCpPi2t0R/7Jlw8n
Qs/yL2s3ds89qnGg9Nu7g8/PbmuRZIq3cpgwYOOTOAx+6zbBLaUSja2q1pfX8qWIJwJaTbwOs484
EvwcqzhsX/SnX8XVCCcvJhUkrbQ5rH5EFwuG+A1afXzPdOq/gXZocflgO2Ry0xxHNx2LqR/VgPyT
7zqI8KjWmi9mY+TKv9rVu2IE8sLQqBGTNgzEvVSm36DbRgcWl1cnWZVgLaYEqZY9gbYNG+kr1mz5
Gk04JJU6Y3tpHCUv4kmmkFSmQuSzctEj2IgyRhU6UNc4IR5zWx8BY1EFxnVvMSzmFdpIpFoVr+lU
wAoyLVTDsO1NyueFNrTg0SiF1OKwXLQxaCZfGIQGjqgeOL6cjBh4sPRIv+A/FZqCd0v3Plh5PMdT
x4cRXz/JErCQ80o99qnu99BpaVl19EM2udk9tCmhoIkEzh2LkrZ6rK4DBT5SjstmJxeVy7VprIS2
7b0siZzUzy0h1XdaUtrj+zAONs+jK5CBdI/TL4Eincc3dG7W03fjpx1dXF8axmaE8GYCT3gHCgXM
0EwMIamOWWok8EbsH4mr7/6YvBMpqBq4Q5IEGdK3xPEb/tpaoZ5WFiSIV7HliLq3+KQUS/mgSJ2P
qpP+5kR6ncKHgaMvqb3/811PsAh3gCWXPDDILj5rCFZIOeIOR2nxIc/Y2W3J7rW9kSUMatjybHL1
xmwg+onmi97L+49BtS6rHxGzr2833VT71z8O/Mg97NusXrlk6CSUTNcn6HUz3MB45dreT3PQaWvJ
x9/eM6252RPO0AkJ4lzWhERVRqUXAE8hbgmnYTvGUcNAPASpr/rt8cvQc1WaID3CYwAusvlsijyr
jQbTGdrrKYlT5D0uigsN/iNATXSA6dc/hB11gP2TDuNopegMhTHHnuSLR72+Y8kxKU1BL3VyGY6t
bSVEmKbpWxsAlR+rNnYbxVWZrbuMFK1uQRMdPJBz2aMt8RGmcErr0CkwFw+jhVp2NvLTJGot7lr2
Q9lF9/TjXK/S5j2di/eAxX0Ps9qJnvym6Ku4jkiw13haQVKNsa/prX987pVQkHk/7QFVYpyNbfLH
nVVYj2uSGOVf4DrewRgj8kRxAoS1x6LG0P02yNDRiUl4GBW3Hgg7zMeiPOVxOo6EqHI6eAVjg+po
aUIizbIsfkVOntj/GP9u+OYnlBy/+yTidi6mnqVBtfdaRX3OI1b2qIbKMZITMnjpiQ5UaK80F00b
F4GbUey9qeh+WTR9MR154mJnin+OmFAj5nFL0zwp45xdDAJ6aO0oCC0McEQL8Z35fSdwtrX5E44i
XzZbTM1BfTeMnGC8hNXjIhz2sbUGGY9Cw4dvvzkIPuC5/STgIHCDzVi8OJhxjDynfJb/F3446ifX
ygOPH2ZYgCIdvZ8dQUh45d65h3vPzVfiAb7cp+jmnvE1v4iEHo7ptAiX24zNGEMl4By5IzobjkGj
w3VlMAbhwDfr7ZNf2MMSxUGNW/tzS21GonC65H6H8BQxaiRKraM61T4XNHhmV/2OX9PFWrF16u9P
+EPuI1/jGfmiN516eTR+gDFralcF9UoJlxC1uZR1pwvH/05tQT8K7GsNAJjisRshqITPmqcuDfeO
X/Hhb2xmtvdenW9iEh23Mg/iTj5/N+/i4VrYQAUCP0m4mjzXbEkDPBjflboWXzsLXDOk/YdT3HLZ
K/Tr0vzc+5UKBsMUKmNEjSzmTfc+EFWbkod8/a6xgBnHCFzHGWbQxZIx9ahIqGVRGuu3HvZQkdLo
oYsCm135WRsRvX06Kgo5/McpHJu1chJ01/Ox4cqowDMqqEB++mIJ/ad1g93JgqM8TCvENqqkbByu
KmlqBBW3cC8zImsi/5ssyBY9gvWzhT7C6kxNYDjEyhdeSz9oqGuwtNN1T2/Nu99B1xsRLcdgWfFF
H2KKMIqDUzIROkcAZU8as44q9d8JE11VE7eDAzzKVFMNFY6TFlM0RcPmovWojAhbJjVKreQVN2dB
jI6HpkYvl4vvBGRzhxmVDpxFqhmaGtTD/BMLYQT/IEt45xLrW5q3eEBQukJdzvUd1QL/TrWr8J+F
KCMGG+Jtgyu2MYcNSYwwP9pj0oFMwReARbItwca3wSWcQQfMSXjaw2RCRGkQdBVqnapHRtAlYkC7
K5ziDlmC8O6WSGkHPv/psveDWE1lxXy4ZVH5BcfiCILgT9Mld8DbXf3dRyMa5L4cvds3uudK/wFx
8nq1+vuvowZjBZUNa/0CSeVnHNYJTRiP50oY6zTz/grgYMR/if7EQ7zEClvftM68uTdcdp6G5Frx
agl5WS+PYoKk8CXoU194/oNreBLwZBaTJnAtZC6JSvF8O092plMeHkZWY9Z2E5WqV1aTY+1Wr81C
Xvo6qUtOJgGA8fWFwUGgQJGuHwYsuR4+Xwjcf9cRULILHTOhBc+mVrnHLi9PvB9wI/sgUIKlfJ6Z
KQbgNu0PkgnU3Fw1YsQqm65wmMYxFl6tRDhtAzl+Pj8sgHf8VCeVuGIt+6i/8WqFOxb4pj4bIyf0
ZCutQvdrc7+AhsYXJ3eqri9UW8jtOckajaZ0jeC2CI0kH4RJ8PhWC0U74l4s/1ZfD4w10mwDjT0S
6clAxayI0bCj1mtunuW71VDasf7esaFQRpsXtaHFn2JlI94QdkZdk0HwqqqPzaoSEynAqh0s6oo/
tDXIm/+YcoSywtPc96SGOlrX8dNUdPA2qMjctnz6VL39fuJV4+e0wKHxIeT+mDscZTEohUSnUy4b
G0gIyIFQ8L9VcDXhtJpESTSc2rFZx09XgStv4gsank9pdKAwZh8CGH40OvDk9mYBtR9qlYFCPAoK
sIsUWCLqtTKKjQdneCtvx21SOuPbCTbM9CkpcIpQvzq15u2Z6UPy5AYRgIvxpM23TqShm+Bmi/lJ
weUbp7eOQh3GLRwMEXbB1E3hMLmu32z/wmuHP+RRfDJJwedfX/4FXYD5mZePfc6Hyr3SygjT2KZG
Yli+YjJ61HVqpE/t7nkpniPQp9ihJm+mbqeSDKGrIB/j9y4rwZhsbo20qgUU52YRxxOPAsG1l6Va
B7j3QJlHR/HjI7KXx2pXb+gbkO2umNG7VSyjasUKYew3PTtqgXw0f7+FIBigFhiRyZFK7xYhjvQ1
IVnaVGMwiWw60PBkX/rVIQLxqTl1VBeK8o+Lodv2qLTD5Chmaif4groi1slxYknJmKHTKOBHwd3j
l909q5aYD3AgOa+53PEWQhK+PReE3gL94C1LqRvwLcyVmdcRMpMSnYDWXVrkaoMi+xEqWf26W9SB
seK/wnJyVvpyF2b8vLOpHsZ6b2e+KoNaz8DQwb0Tl09iI8X3pLWnFn+ouxenBdUGd+us25aEEROL
o1ofpKfyL9JRBjFLcWaFhgwGFWkvw63p/8Lky8tN34aS3f3T1Y19KVtOmxQlLc81d8USmCAXUWzr
qk76Clsn3boBn/ttPZJQ5zs2KKVA7/omYBLaHUyRuVbg8QlBZUh3tDJ4u28JqOD3eR3niyswhu6r
e7s64hpV4xWq9yJwzl0Ytd/RN9yd3WrbOLAFCdVJR22Q8C0mHWMV2P5jZEpoaJhzucg9PHinqXAL
kdE4Pn8kYX7tCM9j0PfzcWtTTgwY5odY5dCqma4W+URKc1XaXCueJwxl5STWNKIxLvtY8sqioHbl
xycuIfrzNHMcdPeM3QbJwV+2XTw8php7PHUBbmHUtM2pmt/uv9lPwyYaRB3H0QTdubh4dSkHkdly
TPGQ4FdsrOD9SHfWxSCvwHkkrLmTKxVWVupJ5BfU1Cf7LGhZny9na8C8e/6FDCB8RTaeloKrqe/r
MJSx4vLhPGqXi+BzrEeGSfYz0n+AOk5Cco9ZJ4HZKbpGSqtBOglSj9Ngevcavgtqf1NyX/jC3WRe
+tT2q0KnRJiTXifdA36BrhiIaK4z+ka0qMkyC0itsQnpyLtWKIfOtlSlRAsYNhEyPvFfRsk9Hs5y
LUYaqp6EXUTU7j9PN6QdgeAG7X+hXke0YB/pBJ5bUJyeQgh/ix1tQ7mMy9ndJY3dHsicoE69W/Ut
dGOxoBfQy6GabFTiLBKrLyGNVCutrIBYyOI0csiL7TgXShBgvDG7OsjqaZs/hELDdaMWDJPIqf7m
IytqOYSij4rbteiUnCY4PVqJgQWjYd30YKni9vWivQ+qckKbLIni7/JwlIhZLs1EWJGrCMeipEPw
J7u7PjKH/jkoyBT5iTmZrc7CjVAhbLfGQjorp51JJhmICIs27xFgewjMkrfYFLle4sS/wSJMH8wG
LWytsQgQqKsEwg9+DE6NCnoSe0lrUOKZpayaw523rzkMmiECYFjw59rxzJHyXcUShSyn+FQhIDLN
oYW9CubVlE3oWqHeyVelk2lATH80jq1iHsTwFh9IHm+Pd6BKhEPgPmuaLCJJsla2QatceyPd7NZy
bIFXwrnKu5E/l6s5qV5hVwbLxU4FrDmFW7bkxZ6i9d+2/gEJCYXv5+ZpOnbDbBDXdiXgJYZDj4QO
woEi7Z7MYOzQXL/ScF4Q34hiIYmnNh2+VKx4zRe/i3akqcfkvH693TPYExGdTR7k2aY5RDbxjeZa
X18+4Iz2Daopw/QR91CwJ22JEPrZwqOdRQuZ7FH9uhVVSFLpO4E+tjOjtF5TIVWwTYJgN+bXa26s
TCgFQVDipfU2EAOOsA/Mq+/CYeua9g85YvfNobQHBzeDVmcMwHwzsH5itwM8OXFSMAuDNFZhJIzZ
L43a4+WdVj6QlnL9ne6gx1g/gRokiWO+WOmzZKCxOgXiBvfkvSM5nRj6j18SI+Y0vXTNpJemElDh
+fKm2EgLt2xPydbtkNHnpv9O5ffwBe1+EQQMwxITO07lRUuPFVGwyr4lOp+34IAqD+QkXJWSej2n
sHOdJ3h46ZO88Yq1uvo2/3hFZWAZfJMwVJo7vRSf73jBT5WAlxDhsEKWz9loC9ee4fIzVJE5y6TE
0L0E9RCgD19+t2YucPImCiNv523HnLymVSDJRSm5GzunJIoIDNyuqYT8G0EHbjiPPBk1nUaazDvZ
plA8QrVE7vFJLSApuXFTlLPRAeAdBnwFI4VoAoJVnOigTEy5z4hpdTvZfm0rD8FnzWpmUE9BKzE6
O8TbKZh44MjS3oRrj1ZfMsI4F7HZCQN4mT+uWozxS7ewMXgxDr8DPZGqUQPc8NG091q2AUMxk9sx
6fDODoF7MkCj8FkKw1mMQGGcUvRjxE0IOcbWF1M80dvIRlVU52/BpUBKa1w733C566th0dUfRB81
ojOxIEgsvGBAlJaMw3o+5GNMA/jcIs2QEZDqTdOA/ffa5nDCCUMYN/HrYokcjBiFGvvNB//RrdFZ
cF2T4gGMBJ0BG7T6MzpCVJ70VQlmWqzEuCikcUrYZB6hpWxz5nNSwCCELhmkUfzQqwCd24e/Ndjt
dADqjZRnWfEl7zlwu3FZziyjo1M7aU9UTYuiXfH23egtzNgHo+T+/aUSUDg53tu3qexKT9dMihin
16Po/ZNrimISL8GyrUcluzuZlE+1Y+1oXE7EH6az+XdY6PpTwj6T8ZUh8LpSoSQ6HITHYIwUHWv6
53V6axon8TzPLSnpCB1Aqc+TzXW3R2euzpxAO4cDkZIJIlQT8ZB+AyyQjGXQKkc0eE8x2YK+1TwA
P0xlZrlVZNdBmikEBnyZLRGQg0khO2hQsRW5zMmcoY4aZvfpY36KmN2Kvp2AojtXc914Ey3bx4ic
/3jCEnWXkEdqfsJwi08M+rXqs87yMa1uyuF+XvrVmuVWdoTk+MJ6nQhSkCBog1EXDjbykijhsmM6
x1pJ+Vos9O7m9EyJZKthFxkgpWBcRV6S/sTMDqitTeZXxRC/ix3HsE5O4Y4u+08SMRv1+kfHdGR0
ogzV+D+zd/jz/BS8ylTbJuqOGjqdO9wzkFUbBbNy+Uuq0tZuQ/Cq746PUvnA4RqUaW8JTwe1h90w
VX34F7TUrTz25nGbzb1I/2KSghcXoF+ys7HvEJ7hDy8mQQkbaVKXOZSnQOkzWc1x/Qae+vBK1MCG
kJ9xtYiqI5hIJccg4OOworuIl8Hc02BmnqcKfI2USWPzp0plo1Lxj5nuNgvG2Dc/DYp+/jxDs4KK
oZImHpALH0TE+bIIdFy8UtZDZICtliTy4B1xvhsNLZAunNC1OlIFvxARtFyTHmvG6wIou5dxnFr2
7pDLj9QUoK5gZwAILCNTcZz3PPiUOwbC3r2JgY7I9dQM1PQOejvQK/ETcrrSDT5/dTsaHFr+Tvi6
f2YIhsHOKwFBqbMs20NlVZrSiSU1sUwxgIc6TueiNk80bXGUGSIrE7352cRzu2qXnshdnLl4FfZK
M06L6q2M7J+xg0V5pepgK9hK7YgJ6EfpzPMK5f+l3dyroXlfpbA97dHgW/+a8jBgqjW2Bl40MB5b
iW3oNerqjRzV7rYHdua/Qbw0k/tbu7mW0gsxw6iItwaDg0jLTQ16KCLbhre6Plk+TCcOWL4FMahh
qzEqhaLZYyZDCInun1wkM64+ScFVwbZ4HlsPBJn7079RQPZ5WjrusgpXZ/lzX9XQx3AgF08o9vgc
SIyf5iPi3Bwfdx28Rzh8EYTzhBH/7wg4Cz/CUTobZBJki2wiLkc7TFJWU7pcT+sYPR+foaF5y7ld
VaQlCFzVGlP6ykLCc9+j9LRsoU4UDQTfiKjWEBO63DZfgKdXq8/OhOWeXAy+YEjnZqFTEWRyZWQR
lPAeasH0Hfsu1Ti1znZCAWYxEU+JSYJ0sT6w42YN8Q4E03ohlI+6zGFLdWYFAmO1FBtTvrUOuAGV
bga1YT0rw+/Um1QjYuZhCBLgOjD8l8k+61TZQfh5W4FNeDfLz0eGaBh4OHIKONjjcjjWbUM/mKAk
0uWxzUJf4Txpwjj/uiEPpQRR3PfUmnD0MiFOcrXDniWgQ/tgTuKFQKFqw/8L4UqAY/y7IdJzHVVX
WVsno0svznVvACNgY9Zbi+9T/we78Tx6OsDU0WGmodVsKQCWX5ZImKF4MGO5KLjnl0lDXRIbLo/3
wPMTSaRJKt+pTG6UJ9Dt9Yy+wFW1pkAiNcZtqZSk6SlNEzn1qtO5wKK8iH3a+Ig+KITmQZcrKSLi
7L9eFfHT7wKoqfr8hHrxi3Jq8kVJ/v7jFhjVfoHXqXU5i+pFnPgXBMeg2zzlM+dJq0b8nYOa2sAa
+MJwGyyqwnB6iahrjesxbW0ycU+eVQlpcpbXeiFYWRtfXSSYjf52v2L5kAyz1sjvj7OMMz91D85L
rHdz3HZcRJCkbXylFhkeECbJYRqDbLk5kuF5hJ07Tpo2mlNr5ub5nmW8ZvELRQiWQtQ91qP2VSwh
PH2JUONUO5/2ji/Yf/uBXlzAZnMLdZ6RcE1DRbTmpWw8871hivRJVPrgjMqJUY2tKFpx8wkS5MFA
GlMVY0gSJC51JI5CGWcGgJCZchnNJBel1idZZEX417/2MhFUwss2D0UO3yJWqyJo7HplHColYjUZ
KHKefetcwGT4csFmOObBOJn8K1acGodKZGdkp3dAoEyIFfyKOETnGdK6fH7vLW9u7JCyaV93fDty
vBPmHE/Rq4YEWVvZwE9GIXqEdXP3vTve6ynh1qbHZSEtOLp77FfKtH7lzQU3upD1Y3kK6qBuYImn
q7Fyc4y+kL96LG7tK/eQ72puPV1xgo3GbOk1hxXBZw5m8gHZp1R+Zcw0Pu/HnU3fOzWCOnAAMOQW
ptVGlOV+SefBc5UvhOiLgSsRt2ynbfzPx0AbLJrCdyLYAUtfQTL29QizYoBeFv20PirFnF8Krs+P
is488hvu6bOScDyd8fpos207rmM4KKZmk9AvPWaLGM8uRQpNE7tubXva/97AkKS2qZKfBG8+T5NX
z41RNdw4ef3o5cHjhUjlnFhT4HLeIaqV5etolJGa8YaKqYUbifmEjrqEubocGYMr8+lJo2z5xoKA
SPDw/a60fP+Bch3xCattZzlWiyTx4y/u1GEgMQlk1eqyQC3rpn23XKLzNcLWKa/bGCd4qH/ozT7N
8qQZjDd30gQWmqkysnAAvGyUzYxMGlzVmCeOZeYgcNyhYwaXQPu+4vt08B/Rpd0TiWvre5+rG1I4
hE0B4ww2wp1QxFL3HqNs+0xh8P2+FUR3JT1VZMZHJQXLt3Go7YqS4Vvz8JMaRmVk8z/W0DqDBmbA
B/eNScZJbLvpPIMcPEyZIZbU8yAAID7LuQUKv7ztIA5LDY65nt04ioNh15c55p6+aty3JA3lZPCj
fVzPezeUGjI8fvVqQ55dathw126LpLg9f4IfJgjClf1Ir/HTG8NE/02LLqdLZRsKp2+T9wdcavC/
w65cnkosxDII6e6s3GFGUpOTtiibDDWa+03LTpTjU24FGiYP2eXvP7SLmF5eQlta0anyBwo7HZLX
oKpnWEKYJTars90x3yvvT/g8YOuDz+/DgxkdAtpR60JYtn8YO7ETz568FFBlhN5lZe04HCu2saS0
CgzQEB3VHdVVlVFQE7nAtXZE92IgJ5jrt9+soQ40zHYCaFlSDLdiJL5wzii187hge+GnZX9e3lqU
iJCe/gZp6FSv0BhYoayCia5sHaPc8ihM0OlNBLo/tkJMSk7VuWL8MVq5tMPk5a7KZy8eBgA1KVtI
d1FLRJKbhjtmGy2WNkjtmxNyGGFQaKjRE6xMwLbIPTXCwIKhyvgEEaiRkHy4oiiMBFFmqw0I6gbd
OBceihkRNGaLHyVP2xxFspmSo4tnmbgqaIc3AP70s9moESr7IOtLZ8roOcEl+NK7LldTKu9nvz1l
sTzsd3J6R914GJYLiKK/RemsGN5FBiVcM4EBnYcwrlUH2LtBh0mb0welr2QGMJ+5510BAubryYrA
Rq2capCAuWPKXdIcWPVAudR4SCdBzCHa5FlonoCqoP30wvnCrlDBXd+f4b5I79BnTGky/xQgZ7YS
HeNJLWe5Tj5s0wajN44kffg9/ZmpDfmKtaR4eDibONKpJ8M68xarxYJ8CFz/KGhPbvreq/9Z4Cru
GjTef3eWWfdMmRKfxQvGb/9kBTphX7jS55i5XpmA8oA6sR+XrXoNZw5I81dFCUe8WA+8lNUCNxNP
Ci9PW0gRvDNp7wJCP2F+hlJKJA5NSRWIT1Sby/ubEdc5oBk7D4DsHSbIWkATFaC5t53dPiDCGjTx
wfZlkb5WW4g5MvrAYvbRoNif4etUwmIkeuQYbRi6zozuPW8Oz+eOgOrI2mcgYXOPvP4/qLakWm2U
bU/sX+V6IqaDG5maKojWpLaNn1nRZcbO3r15L+FYwLK1kGw1ToupcZ+slZ8NJSZ6lpT4F87xxkoQ
XcZtmp6ihASdhU68NSR3zqWjNUB3IycJ76LRO07ww8Nu1WmLYcN9YpjO1fuEjcIOAEkd89HOom8A
QkjiWlIP+e630scVfYf1ulo9xt0EegxwCyKdRxzEtwWCIqvW5jya88OBSSCjRfv9koebJRBvuq6p
jMJSjvzlyq11mSlAULvbRfK/Q/2/0kYjjnBgebwS/c8GMBJHL/F9ndyCvfuUuzxdpZz2AAJyD+X6
s4kOLDS1kT26cnS9U7uSMtjs4Z5hWI7aTISKABZLs1A/oW2HGrsH1q9RttjUPVqESXWk5VSEgFLi
66pBPFJRt5BiTuYtZS3ySf4SMof5jYNmiCEldKXRAzQXt9E5LCqq8al/9uLI4IJRnrNhZYbYdaEC
+EPpGI9K0FS9rSExZ9wvntkcd7kJArB5ijvX1V9gU4od0wD1qs/P4qGY0VKWVSYdfiEilOEtE1Da
6vn+T5a3aQgQIQSMA2+d4s5N8xzYuzbFyMjAqjOE0Wye9dnx11laTBVILNYeHt2Aupj09RJFaDJr
bvPMvqrXRsOh648o9YeozOSjmtB/drfqbOhh5lrzC9IJjpn8F4FcQdGOArYaIfFmDwUjR4HD1jcu
xtQ/R9xf+NZHtzqzLLTD3uQQBRZ4Ll8iLx2cYOBOU45E8yED3SlyDCPeT6JGjyIG4XoqcI2dgXl5
rINMJ7tTqFCEoXptoU0RILf2kugDRpmjeM1B4oBwngZm/2iLK9ty2SJ1w/nBJVTpQMi/JSibWq7z
7RI5+pHgCxMGz9LfUr7ydFfMfdsbzQJkWEbj2Nw7fpsgTqlpQPhzGPHEuVbwY9JRO9xgNjNgmInO
px+lhItB05KUCrNjg3iU9al1cPaHVf23MmYjDTuDqrxPtYzyvkdrpp1C2YMuXO5nLzAzyvOv4Kli
N/SAUw+myRw8fgSvrKVdtU6AQY718laKDqeJ0O5J9Iieqy6hjnF6zkufNC8PKHbIfhMCBveLab2h
yIRoigm4AghPuzMATr7JwdpTXhHD0J9ozo7oGbhXemgYwwWCYQ8l0zURiUrvSGj8dvGBIT5VVtB9
1A1OC0Dfp9ELvfk6NjAIeIzY+VpoqiiH3WiVVtR9xNCCjsbW5JMIDk6n+wHuxeI8in55IS9QQefi
dk2/mpSI+qbDKSbxPp6dFm5ro38MSsZFiljyI3t/mCHNIbAblr0j7Gu++gUndNoSW5BM6xdVgxKm
YdwriikXC1oa3RjARkqw/Lo7CXVDBOXGbm6vCheSTBjHKBZFh/9LPhZxo5/f92+Grf0WM//DsEBL
AzhGrPDl1N50jxcccz3nK+HlYIwJQsG0pOK4oS9cvQ4kDpxDkD2c7QGa+ntJLCpxBI28HYZUyZ0k
E7ZT5e7xqG9lY0HjhIEf7b6nLs/tgLGzWX0ZCM8SgWs8XT/7yLNxL8rKwjw4JO/By8J8ySx3BDSp
a+UoG1qBPFOTk5+bJIt3p1cw2odwxbsB8X0fOszB3vofuLaNbBN5CWPWlQM464yRUpDni1UKbSVa
WbW4px5AhWwxxDHPJQoQtIxC9A5KvMxgdIEwB4s1NGvi+fBuOJ5/iUT4F/oAlfRe8UEy9yZA26mn
Wxe++L5by2IfzG1mIVuY+TtJdWLlkynBIGeJhZO1ahVRY4U4SoDTpKNNJpzl4xMdzCcpK9zcDmsx
XAHkgW20BM0blXUGvr+o3EGFGw8GExuWgPYdeDAQHXRme5+iznv8Ltt00yZhJt5MW73/iiHrYdea
dHG1UHCO4WaWQNjs0j7jym3XZtG8pnqSfGYQp3e0IqSn7w1gRj2DxmAqyxEe9yygJLCYGg2Yo0NP
pvN9MudWAyDLSsKeuHTZJsA5pPCIyD7vr+74EkZ/e7R8jCIkzX93Ez18kqAy8hMYQmDmo9MZ7c+q
6vWz5pmcHkXajo+oa5cF0L3jS/kQQidekLVcNQfEG51ZqmSlUCZop7GomQPtTRQMYqvBe5vwbVW7
O0ByckTVmf4Z90SXcI9c4BkxPZD2B1Ke5+psZeUVpzFnbN1gfSI6UIAl7XZFLrEPFAr7MOPFa2MK
3HM1Lf2yGvkSsh/JLLeVM/GQLPqbDMCtoooxa+3dhMt3XNFE5hjEQdBFylBhB8EbQw0Yg8Ridxw2
8ZOTmxf0pACu9YtRIyj0VI9GZ1jCSYExZdAA34FCTxe8b9XbC5XnS9fTIwq3PEoPKUH0fY9G1pGZ
3uAHgBc9gP1L/RxDkXgBZh1mh3I5BcE8+AD2qpkHpp9R0Y++sNPdkpcO/4Ui4Etr07I06agtS99d
X8FwYyvn6eXzjLqAdrn03bojucLMKthxdzRYImTzCN6ej3s6RXPRUE6H1qpVba4LYh94Gn70OgM6
jVDwxjmgeCAhBmrVviO5Au+FxwpBFQFYSg7OQS2DKJzlHwny87SZmT+qPRjRq24jisrN8XD+g46i
l1tj0AukDglCgBw3ItuKrJpm4aItAHfQq+nHxIDX14PdgMnB4Yu53rzLO3ebLksobaE2Ze+NkDjn
gESt1XDTKA1wzNCTdsFYVqpfQf7wOogV3LtaHIpTije7WPvQ53Q0YIdn0ofX1ZZeiWVT4cNuKG1h
r1oFrW9qv2rJWDTgpTn5j9KIjwgkbKkGFqlpEK5Pjg6xrKvz5P9vUlCt1rpXALHgb597cXyNB0Id
uuNpNd6iPAq6kM00uN9K43fBTnaC1AVAjZMHazpaLpfPvxx7CPqtGp1WixY5l41QKE/Eh+UO6C0a
QgBxEEqFPTOjzFcMITScUF4WZdyCGiAozemx2jL0uCW1r0okE5eIg11Qzjd2Wj4UVqR3G50KK2Ec
Np/ZRJKfOz7qDoM0copWGN9XdwuXOdpjRiVcG/ZSq3x63Lytjf6htHzeL/pVnbwBS4aVVZ/Ruzdc
QBhkJaS6CWe1t2eOagyXLfChyuOwuvrLzZu2cO14aOfGDMzCRWYkmySbpfzU3t9E9Uh35Fzm+ZTK
/Gqfype+/muSacWhehqUilSQyItjij6b40iArZSAP6s/CpW/XWMBcGk98n5YEZucgm1DWppny3Oq
p4G4cRFccNGF5PT9H1UFjA49rB3OmSvkOQegP7/A8eaWAIHE1umbRW5ba0mhpykFKrIv4U6uHaF0
RDSjusFHlbsWQ9es+eGKKfwBQUgQHSiOJn+lgFKjOehhxg2b4XgV9UF84T+yxMB5GzN/A1L4t3Rg
v0P2lNePJhapxHQmoWQX+eGtJ1Pt1Qb7pqNDyL1BHJbcBUwp0xJZufRS2/eLcDCiLXKFZESbrEsC
QIPW97g9rycWn2AT/Svoq+WEWYrtRhsBCV+aK1Dfa/7u//iX58A3Oztvl4yQaeXSVF9BwB/5/ZGk
WoSEAce/cpFXyHomhFyjl6RQbRbIDGFjU9QbJnkb2IOE4BiATQrraVnkY/B8dLYTJ6L/1Vo/3K5Q
GEX4UDC0idm3woCDTO6D88Sem5BGeP8L78m8XWqJkAgSA4XCev2WXbV3jSWLlsnMJx86ZEvmxg9O
s9G6uP/UJU8ZMs4QN0VgWCWwGfkhfqSl0673jx9GFJm9DPUIbV0tmTAiQK4ZSn0l08zADmQ15phm
9hSdotw1kyV46bancEYE+keyvmyz8jsELNnHXKnTBwhc2ck7SuogTMHcptgaZhEVeAUp94tLPLeV
0YDBZKhWwOWKFlGR6gsFwg/vel9yBQt6FuhfcU2D9ShWjpCg3lyjPkmw2Hh2zzyp+28DUy6S0ccJ
rY98aOcL+E+eBy+D1lx/ZeY4J2SBBxHAw2xP0crySn88N5uT53UiDCYZ9if4Z4ZNVRvqaDQ23mep
FRuewlSmlSJt8OuA7EvvynU+MZlVYP7Km0Q0eAr5/bNCukliszt+pA2BAw+FVWos/eL0un88fBBr
bQqnXhqFfkOCFnHOuqvLMNdEvnh5N8WShVyn/LCJZndB1zg8xzrcE3wZLrrDvTPenheLtd1fTTkC
YWDxJO3iMUfMAxHlQqwgxeT16e3L4bryalcwt/QXyT39wNGMiQEBC2seEhNkWJnDbC0j17jX3/e+
r5Vq6BvnxChKaxZ9siIcmow++7ZsqHbo86N5kNmokXnR37Ln1LceH8FFj6PvkFLEEXXRX486m/DG
fBS57EpsHoGz+CG8y1fHJIbcOy1J00PHcOyX5L2MbG8Nxxpe0Kj4S6hCuYeHXPfrQwdkM7aTHvCW
Yw0C6bh3EATmZOXuAl56d8gJhzwbnXkmELSyuehYcu1/M8UW0V+XjeVcF8NJ7lhFv/aoulzU4Dob
aimsGXLZ/gxZcgwNWfLCCPYXlTGFCsM5wsmOemAaxfsiOYOryTV53ldhamxy1jlItF/pX2xIlUvB
F1s6Xg+kBuNXTxHgYRr+qWIn1AB+cj2VAj+uSw7WrfcxFJXpiZxcUdL7hCbTdoPs3hZeGUKog87+
A3UWcF9rxb1+i4fSZDi/eN2hS2D3LI5aWdZXtrnvSeMKSSDY56NoD4igblKgD+hhVtL13x/U23Zq
lhfp8jGxDgZ2uG6BGBpCnd6K+GeHaAlO9XsNbRJs/49z6dVU8LxvP1JQYS8U7VVmSBAr4ORp737R
7Jlgp11AzJMxeZfJCrawOULmPEl4qLGPBWxBlxloKCX1WIz7WFZOiQTn5q0XPcLby/+TpZIb8n0/
8Y3GKoUNER8ljPOtY7agmSNQCDdVsQyFKXZUPDr36S45BopBZ5mGcLkLuWR2Y8KgM+mOigJZOErA
4chxMJaFrJ6pxrDbABwyB8ekhCSxaDEugTPVnEZN/rwTJF0xnB6ISyjDZbiebVuChwYt14zqScH2
8R54AJ8JNkbtWUKV3R999Bs6tAqH8+HrOSNwzG4svqRDndWbKTR6+eOCfj5yrScv2qvIiRsNymWc
0uQcgNx2nB3OX7/6VqOzwDCH3v0fAFy4coZP/dOgj9uB+qdQIsuONz34WVvWOhkwpJx7kOR7QMRu
fY1NWQf+qnV7OyMg8fV7oJoiVUZCf9AGMFicc5ZD6I8PJKpdkR0SIgvlcSM2+m58sm63WEeYbRlK
TPMz0CfSvOxhxt1CqRoajN7r7oyHs1dcBdNtSPtLgBlWnBBraTHx6vYAHxwZ6161fvlcKF/fsQ6e
MX+d+V6qG1P/UZnETqvu3PW4IOp85+vcLqiMhE5Up8XXz+3k+H/+lzMFJ2tGOcQmdVrFQ0GlmuY6
dSNy2wLIZEB1ejd7+Z+zUjmFNi+3XY6LDpFb6C40BJBjfLQZkoW7wILegFYq1wJR6c/QVeUSWVra
NXdBAkxuJ6QkId1kwylxEINMD2uTJpThQrWVLkdeHPLML5j9MDm5ow8DjpQQW04RZ823PM6xTKsS
fNFBiq/QY8GhuPCy2kHDwe0d1gdXRjiRiqzVMSRtGstAhR38p/6JLNQLPx5EUNi8gPPlTOv4e9Rs
iQxgQ2i+/gpaEb2T77F9jYygFe/S2XLtMVSblSzM3BaxeLyqTylhtDQf8hJv7SWc2NTzS0SNS6YE
aZDpckDT6XuV4ASQUq6r7a6548lqOtAdpwUwHcuv7AoPxbCBCsJR08HkmT9UyI7D7YKIUtQyqLrF
ErpT9ogVrHsl6Y4WEkgOGsbEV8vJk3i1CCjf5lI0jKminI4ROy+5Iq9S8G8HBxaX86FOAPaZPQBf
p13ac8BfTa10KUX7tpS2UUDCGhA5ZMP3jlph98OJRWbMcAZvYX7ukdju/acLC3F7ceuj0fMz8ilR
CAB81qZ8dc+Jf2rro59ZJr3jzNkDXl4iu6seu+ukor9qrej5WbDc2lFJJzL6gCslrdq+z2LK2QJK
KmBJyzfXPd2+2H+ViNcB+k8lABc02eff+awW3i9VgfeZifUlz/IY1pIDStiQ8zLei+VMSsVvXMZT
Dn7rtojOCIVU/b/Vr0xlI2vClYAf+CWljIITf3BsHzCWzsrhKjKfNAaDbNTtbCKu8VUoa2e4cQk8
QHr5v35m4raNFSaoQVapRIRqj67x9Eqr4PItCmtU1XR9P3451Ib5wtD24edGDFmKZNA26Kwv4KoK
e0Jhes2lmjBqlVKiKmWbmXvNzr9LuJ93KhV9GSLVEsv1QaHGLbd/dHv1npcfFtkCFZWMkVv40Dj6
wQgmRM3x5xMrBMnu1B+0+Hs3BK+bMChK6pjn9364gRUg3BlGWHEPfFr+a2gjxVDTWHCRLQB2zizf
yZHCFbeKHSHOwfLBavGeUG7oLnLC/gXwEXAlg77Jp6pvNx59O1gpKWibZTnZBFIBeRwwI1VhIC6c
Sqw2+rVSmi5+zzjsI/lNTcqbE0lQ+q/VBu0u4CyHoeHpfntAphjsoO98wjsDsS7mTGP/JX47DGbp
kOh1zx6+cQ3NJRHAgZpl0ZXXiXUS9fUkPAfsrqGgqlI06NalZgJgmw6dYcWM78/r5u+RspciJyMI
cLAMWjyd3+/n0jdFE8W300e6asrs09iEJVuzFI6ZQccdbVNrpCwEOEq1razJ/7GKLudCuXZi8fQI
scoU0cLgewE8FfmSvhEgfeM8AXV2KZbV7RggO57IPfLx0gy4fHBOXRKnTTSFAbqlbQZuFBi63flm
WsZE/ANDSkomNxnpshP29U+APm1QgqXtPS6ulvOUuS4vLM1SaYppPtEFs0hheteiCBt0qWLRfRSy
ge14jML4K7Gik5WOfjwsFVj8T5BaORABtpldJnDJKPgXsRkKDM37Ka6uYy/D3v9bh0V2DQxTqFRX
u469DiQezp2UuRydUJa7YROcWOenR3v6GboEeXWhyME+iTFywlOqVPSQFl4IQuXp4ut+e3pFuigx
z0skPekqZAxdywnB2wP3db3Oalq85V5r2wJlMbROE/R3IPmxoo2h3fNLIRK0MIuzi6cb1Umlwi22
zLoFgeIpIadqSTZbuqB6tSvhpO7r80u692sXt+530BWRf1KDYVfx0sThRy4g3nHXE324w3P3BCPE
2CNFYHEJIEXhAF1CoTvcD9UtgVO65U6m3/Q5GykkFg/pp84Ev56PyUIn1sWmhqouFCZv95nLaZ79
UmT1jIug736tQsj2ky0yGyAC0HIf5WUZbPh3DH6PWawFpJiOoazAfl0U72mfnHnCz8io3gSiruC3
Jw/30wAZmxVF3+BqjQOALzbeGAkwuZ6Qv7eUWhL1j+IMEUVENhmfr89n8RK9QbXKCLTJNOZc7fHC
qg4VIKVr2qNWCMlSBFwGhLZ9mppRjBt6b/lPA29oinFMFFtMBKlZCSvuWEM2h5yRi2Mv8ThoN/9l
KQEgVWlHfAE1m5RlDcNDKpbeRz7qR6NAgjp1XVcXlAIKRxjhD6zCk1aFHNXDQCIk98QoiqZN5Ae5
uvusyLfO5qEADK08+u9tfiwRtRRKq205+K7rPRkmRGnWIgcwMOK0jviSTDC/A0Ni6f6kWOVYCFuH
nF5zZlj2rjF2qFH0h7wZNuv/mZg4hNGwhh0aPa5iky6T5JbKf2C6SS/TZdT7BZQq/xy7TqMu5xBS
AymoieJLWojdNXHJpC4CA4M+YeEgQyAcoP02NpS7wd96kxcW3EcDwBxEuG/dzjDdo7b4bVEkG1K2
YKiUwA9HtvtFlLB6RKoyKzl2JKFSFNm8Z0Itk9RK2u3gjDurq59TgFs2h5s38movhr6X9URD/xmx
eHSS0LWU1vOjC2gL6J3DmXhimufqfjViJNFTdbRqiHPcUvcY30p/9QxBUbykRAJ4RYNLwLapi3FH
nXK6MXqiN60qgMT9yJ8VAqdtBnPjvOxGvHJhiXBT7yy+y05DxhuvfbOV+K7GCHyX2a06SmTU3k3L
Nn6QFQKz76xIawrZsy+SO4px5wl6wEpD091EYf5NQ+IL2yH2tGJsLf0uNa6A9MQA3zSYAirvHwev
NbpME3rYCZVvaC5xogrLTc9pFspoGZs0soH7VdfXe6VnG7NB2isGj7Mq0zQNViD5KZxRGNUlsNzk
p0Wy2qO9ZzzZ5ZIQDD7hukUQM/jeaeHXWlpaE1CfXReYG55QvE04fdxUXy5si7ZS6IZQEyWWvkza
XX73qLJKLeXSKyMNFZSbUjjVt/QZJ7RKBSz/30UIROFY6oCg2G8qFc7hAwSeHp9O358L9is1E04B
BNZzWRUQ/ZfpUM+R3o7PJQL77eFq78SWKhsmPyKLU0yEww+897NysAyPw9g0nsd8WFc6TPlLY9FS
lpIsavV9n6yjeiVdWMlrOd/R957Z6KQiw2oY9ylS5YoZb3GuW6SL0jN/l32cQj1O6FjWGU+OFqGd
aoQ8Zr2tqxCZs7G6hZ3Vqdb8ZC+ojnX54h9oN8u2zBqlG6khaBZRRWbAbfPbvPpuH9qrtq9XVKaM
fs2P2agfwUg7gmD/hzTQ8iOCjvzrqR9ub9c099/PJeKTXtK27PccvJBKub0SV38sTi0jFlA5JGGG
TjQqD+9rHfNBwiS8QUkKNSD2yHBbVW84sY5/hgxGZx4SKdpxEU425xqBQZLDG4X9H/iSRfywHAgj
Ij8cd38xKULrak0kAm647fH0p4bkgDvSnNBUOH3ZWTLCjRv7edFLgAhAmBc4ev4/jTdU/+utFDEf
heOiy6SG4TR3KJcb6HRHhD3COIVXWCNXOVXNbpacmUza+G+JErZp4JOsDHW9LLiseZjeLlNG/46m
c8G1iN3vcqsoFCJz0OMF3Gfn7dVaRlHdOgnfqwsX94ZqI/0b1dSrp3BqiPvasfi/DVHK0FqP/78V
u2OOIohKAK0b4pov+xMjJ/oWouCTyduAnG2WTuPlU3nwlf2+L6r+NdNaET98p8HwFEwQWEjf1LXB
rQZboC2hExuHGPfsVvRiwo9f7pbGmqJv3D4GiFqjNOVYjchE7DLVFITS9y3kc6rGiKiDIDV9q7Nx
0t5k7laHXKtCwlfjhrPmbfDs/7A5xBGk5GJLtlVXfZQCgjUMDXGZO3OObRZ4gNBO1t5wkBgvob/a
X3b9+gctvUOzwPiJVQzRTS/vTQswSfpT5RtbUPk4akEGB5ZG15G3556CKx3F4rcjdOJMPyDOaedl
5dHi4cJR75Pfu5bSx1YMvtW8YJeAhAEAuFBD/qfB/ZlQ10W8Lm0m/0CaYP/xBp93iw0jQlR1IQvp
LIQg0KIIdDypDIBMRo3sCL/HhXT2AQtW8FlRQRlHLl8Urh39ZMXA6QNbYNs0JEQHS7pmY56mAmSF
d6Hw4d9lgyK3Oru/LrzEYwSkDVZ5be9gYL4Bucg4cIloisz7ookuBFtTwYOnDq1Wjr4oSPCPdoJ6
7fLGc+eU10qCJK3nZ5GYdipiE+HxJyDM0rwkO6qpt5gyf90nHRVj4cxfG7LNbd4BH91Qy9Fw7BsE
7E9BuSEdspvF78gO8zx6SslF9sh+fD0TGMGmCmQQRCVb2WR3LQOfwXWIDrOBuccjHpYScsKeT9nz
cbhdYa/NVj3m4pjmt4Q42DnR2xguSPNCGyOQmYrnRpma2Lu8EIvgaiK0kXCJwI4ow6nl/gxOZ4D0
am5UNEQrH5rnCQ20CNsPj2vbuNxmYJIfgFSXDG/GGjjJaZNonIcmY4CckR+02jz2/kzVKgvFFFWe
Ut3S+iMRqsw5O84kVfienEQ5BgnKvKsowEXPXRMpOlX5rxV4FWwUNlGMiG9e8HiOG1Em3Q77wsck
QKu2z7HleszuqfrVebCpj1k1d9D5fEjFxf4tT/9cesoqY15b4i5G/3jFhcXlA+jHOoJnprUSatNJ
2DSAwxXn0Bj7mzg4hVtkcgdzmKkM6T/yp+E66DbQCDRQWQMKmqeVw/KV7uUgQ5D9Lopql+hmmixW
kveXK0d7Bq/o4RqGO5nLXgcQA9xtuR7IXXMe+bvpYBN6imOf36BgVfpByUzfQe6/WYAFI6METGce
g5etBaQYigCz0gb7fyJX1J2NFe0xZXPgep5c4D93jck821GZqD0gHB1y2MC1pFQ8CegtyAFAk0dC
FrV8FdiCfLeb5aCinfqkcGjvsBnWpO4noDQCPWYuAv8d+eqaIZtIzpvQatqiZ7CIiMf69lfhQZ7V
LxnVaqavrUdaUu9xA0Dksbl2Gmlo84efy1XIV9A/wpM9ge3/kqXSrL+JuNjiS2dR5J6+pZZurDQl
QFyuLXHlHEUMMVOs36F+R/WwD72BXyPQaLcWR6/vbVPmUqyyIVFdcMkKNc95NL/JAQONuimDxfJj
UT3paatdgVkf6ZIgTSNGRS6LpMR5tK/PMVPRXsM6oivHNdtv2p/vNUS3L4OYtbSZJBdHevGRgqO1
SzUmZpW2mdCz2g1q1gBS4d9f4A/1KOJPG/G6wdMQ0oRCNPmqfISCJG+vhw+kJ1lxhg+Gn7hNz7Xp
Kd7N7JS+1mStzYwk6oXuF9bQ1/1IG2o3rnEetV6LFLM5lV0URSwQ+cDP99MOnFAJNWNifZKjpFla
fjaLt8AuAIPvK2yOoJ+7h53PJcOvf+SkCJs3oz/ri1ye8IDn2IOSyQ4wtqWOV2QzS9jgVL4v6v5F
rqFB/8/CMq2Y/LnjUvB5CqgBEi9UmmSzURZc0rggQ8GBjxJn28GEBGB50qRD6xN/AAuuxE4HNWHg
YbuwgeZOaS5VW2gL3zi+TVmL2pHBzzgPhUO6sZNGo+oUYNnV1F4YwWGj5oSvwMBT7Z0qnYhm9+Pz
iDf41eQhilinJnlNTOB1SBYPsYQ0b/mNrg2RCBhPHLz125AyR5CWvtGl3pO2yihPpA/aYt4UiqwY
+U14X70gaSmwMtFQApvMDIzYI3QOcZFqbIwpM8SPkEuU2vB9FpjeQHy5rUEMeL27cBKo0NrFSVsO
aLaod4krLL4DkQz8nx8NWF++KWIU03y/lNU8EMOhsFAv+tHiSZfRPnJxgyI/ZgDUBWn5SB+uIu0C
qX/imtW4JIJMnFDp5QwcuNNkYYfpDkQbQB+t4bzxfWAGRvq/b7HmSuAG4WVClGtYZcK0Mb2TJIiR
7tetpcMscICUNJ2WZ63yfTvIydu0WYO03Ynt7OUkT+dbC3FsZLxPUciITFmkAntK+4lcUV8Vtpyc
awOHYp48vNdomzwHBKO1M/PaJMEuOF1TyN1unDrWJr/zCgbJt4350oCPWWv+fg+ifso6XPc5r3ZL
y7qCJEkhsoZr12jaXktHW8O0GZQxxeiEw5A9L71kn1TJr++gUj4LkcLuhg6ANm6ucgc0LPGGspai
6TkW5tJK5ecYXMLDiZl9IsxVzjvRE0SkXmXbA8FPelJCpsEfTSFD++QCKiau6erMMynWH+X4O5t8
HDxgrgNxFsntWAXMjjEVfDj2aaxhTuUQFur3zAp+QrCR/uaeV67PjRmkverGrdhzRxXuOMx9e4hu
I0xNamgLcaG810lDU55xtWPe/45wRdhxpiHzhHyuTVuWraWtcMKWzy/9AvkVW/xX54POY1ljCpRb
1hBmGldg5T8YfqtLoS6rjawXEJhcpdJ0DxW27xFYfboTQDJM7XW33vk3AZSOGGByhZOwd5fwtINu
vufsqFyYwMJ67zzHt0zBELZZKB8tnAT9IrfDvoq5VZkvVkK8+DU7zVY2ODO7YMmSu00G7uDKd5A7
eyHktDqLwhT4iDyexrRNJwEAF7bngt6rdSPjuXQkhqlP3IfQ0uxE5ryQJKou/G7gVfswZvK8vr+m
FHw1j6r4qUid64QD9Xe5Q3EcI5Lb+TBg8FjeMi/B4juTsz19Fejcz/SDbVSh33md2bctI+ZcjNMn
PpE0aZg8hOeCvkq7fCAYFj5M82EFNJ+EjFPp/ztlSdM8XOftp6Q/tUaUDsCQgzE+twKwfIkP0Po8
Me80T3t1rAGfUQZxlepG671X01ZprOqyxw8+BS8jTOxmyT9BvttfiXLybt5mMBP0MQCgBTAYH93R
PCU14RcV64LbE0dkSUxCBrcY82ZldtXZ/qBANM01fP60w1TsE+dbznSxkiFhx88ngmly3gRB/vEw
jm3TRMPz2ULlNyxBBblNpycXzquEwRCs7UOu0KITP2/P7hB/FKQZv1Yn565uPQClIXvokaKMkkcv
X/rMe1Q+Xu+n3lXh+UsQ6ojOVAj1t+Dhk9QmhSq+v+Z7DCShAMEgiat5R8nLSOoGRPqtQ4ST0sxP
y8K5VOttVpBTd86xTI9PHL7cmwluW28Hi4sW2aEo/zPc954qL4U/nK5CmwLFHe1/pLSrXj1/PBAl
ClP0wzDo37VqvdwqHy/+bGMS/wVpLJfU583xJOBb7nyeErPTnlJeZEffsNhrAcZK78t9S/ebJWFX
out6bKFg3fi0eLclqxOSMFsnyKWL4+rXYnq4N/9OSpoOAB0Fs1DMoyGgt08JfU97bCWfcIpYZR0t
ciV06w4+tB/COdUgm/sUGDdBnsKkzOaysMDefyxdoCL/07OTdaJmI7snfelaEiBA/+y0c9ceFqMg
JxOuPYbSRkvsBVfMqDBOFw8EUNLPnyqJIfdyJo/cM7Z+0OWiX/WQdk09EC5D/Ym0f3TYhSAJz3eO
vot0bGFD3GINRjDchAu7S9PbOpWijjmm80yL35lv0XU7fn4T/s4XAYuIixmdjsmo+8TkKb8mB641
+0FR2lyJe79+jHCkNLXKg20Jqit1fIE+NmSZJ+47tDbUKtC0U3vuye9sxZp9EnAEsqQA3grnpYnh
Xi0oCjoBxGHYNBv93DoyPRrZaokkm5JwmY6RFvqiHaI2PVCdAc9Cfn77+qoo5k1cUpyxikV/uBa2
8I03Ka5sOJsKGJ+3w8/fgqbB3Rr1KAEB6uO4+/INV6rw15nMki6RBaW8IaxiT4NiXHsETs9+Mw/6
CvA8Pc9Ek2kXFFSvVV9pnGJaDyRYIFy9hZrTrA8l6Vtmm8Coo9+4mjbfknsFPFL9taeZY1Js+5Xh
1ORCefxdwO9tWOwwMkuJg4/HpcDeE+BVHjuTRDqkas2teJgJOnbYlyUJuib27HPHHCnbvwDymuxb
2KDgDzkZ4wdsZsJtu8uxTK3B0027oORN5Pe4ioNu2pf+5tmtslCZPL3h5pos5bBOMAA1G5a3xn2g
a4eot/yXVoIJLWif9NTFHQuYEppgJ5SaN5fEfovumYxZE3/BzdzftiKy+6Porq7dt6Cze5SNuc4A
rVWFiW1e69gtKLhgmaXhb/zcGazunFjC+KGYojN+UTcsmGT5q9qzXl6+u38ibMpxIYhFMcmZaWhF
ENTIMZ68aKIRHQ9DXYodggPzcHpj4XUyoXOJIsTwu1sQUPmTvAXEyzwYm+V0WvWDb+uepjTkfnws
VAm29Sf7nQv0+PRuCE/epTSulTdVAju4XWerccTNSIQGX506RAAc9mLWAuw+//TD8M1Vb5FgwGIq
pbY0EL9FtHjAOWTwFJn9VBVXa/q4RHsPxQE+Ph5bipyn6d34CIUMPFvtNlbu1bH0+3YYEOvOFUNL
KvT9BIRA2lLdkmi3S6p5knHGLJEVdLe8HWER68DfSiYDd3g6zf/nY17p9DG5iwBgDbGJQV0CViEj
EZtmUnjRoK2XLf3AoKzWoS1fUsm2AkxtFwtS+BJoft33i+WZNr+OPJqfd5YbiH0Cr9cokB8BU8UW
lghJk0Za7NB6asrj0BQTezuW3wnFpxTsMcU25vsvDsObH6rfu8WschQJhmDW5ncJ2PeHrPuh3+yt
sSb+VzLr5BIwsEwlhUZg5n3ymECPL6NeyEdEBvVNTODj9noGYQfd7ACPkGFOutwE4TA4kTwXEOU5
K6y5wGLCezy3Uf6Jns6k6Y1ExYlTD5RyGzorHSUozMUcbkfx5zD2jhvpQp6Ch2RBn2MRFo6Gd8+L
vIUUWVOp1Hr70fGMlIJa6ELthVXENbbkdufziTF5C2EDzeRbH26OjDRtSYYJG0VAlU/fiV3xI/XJ
AK6EEFjq1LHJs6YHqO7UWwms+51uikGqJIRtuaRKS4ZhQC/zOZE0HgebQbuLhJJ6vNBF5B6hqTWQ
pyOkeChsWMKlTlBU/4JUIqboES9NufYSsShVV/ixbcYGsRODi7jqTRaWofzEk7rGYgtgnJYhbeGR
E/AqrgD96bty2OgH8jyFnz+FbU4Gyq7LeVfLQoCsznRkKzVbj7c6sgQx6uDszJBhO/yhdh26RaCj
nyscg9fqP2Eu6GJa5wkY1eyn/U4FvWHtkrTnA713K+kO4hyhU/QjWM0yoJHmUgiFgZBu8Dksb3c2
wezX8COoF78OW8nxw4sKe5H2dS6qK742bkgHuYNPaYeBFTcjQoLBpdotBzFe+HvnnB4pEoWkfuFX
IxIoj2vBVAOZpY0maqpjaF8afziKYXVu6FgmjoMAk17vYVqsUfrmvMWdph6x+1fk+Bh3rBVKO2WY
Bs/t9WdHL4d88UZSna1alb4mySoWLYM4hLj6plecz0Y4TMvLYsmAxkJH3SHF2ueYJgXnBK1Bxd/o
9JrMlHlkV+8N/lHTO94Nt1DrPhD6gGm1i0W8oQMW3P+nSAmwRsewk7bpowiozeoYVGzvp0QO2iFZ
yZ1TLPfFhMbulhGbDUMSQ3KmxuFZQWyvmdC34blxGwpsrsLsK9FmLwhIxScfiPo5+RtfuNBMP1mj
i4y0kUkbYYtqGQ7b+muoxCeXxV9K6Ahr41+WossFrhAkPVtxpVACBXDZPF1qTa5n1tQmyPT2BGZK
BOc1CG2vWLZer3/N4d7e8cGiX5/lbjhyaDvsTfLk/AW0fMdRi0EKUGY3JTREJrODRc1Dzf6fCgYS
yk50v83JWZHqIWYwliOJmOc0mIkgQ4T8C0aC0mtc+NFS1f24rz7EJfzboUhA9Q59x4xgm8Ac/ZZq
9Njj5x9ryexWO302HjyMhvI5JYYQ+B7z7a72t1zXVH5/A7t9QHVZyn+hToV0qrVcNz+NI31tzkGm
a501hU7U5OzTFUnZ3+btXVMXBEVLiYFK5uvn5PwGkxwoQ3NEZ5ZDWsD6umkEnBcPQe6jqOtMiBNI
YOBIgkuiTc7SOmg1WMBO1pgZbBD/yKy8V10HPWgF4+Fa5zQQJhwEGidgz+sOj8y98ODoZ2ORSw3v
/5R4gqjn2h0q8gfGpYFUvRohW/OQtbcUgeKFoHR8sKm/uEeyrL6c4i1WXmkcQCiAooIwPsYBhZ2Z
Nm8pFXBrBZdPO1RbQmf3IJ0KPk55rVOIWTDLxHLi2CwNFwFBQQ/zFzn5aBXJ9Xf7enYlxaMEj6Jt
RYO5AUrFQBC6JNbIs8L9eS92+U1WXCUi5fzmGX1I3gFlP1ohoguXgZXUYVe0mkpJ9BEPZN4zUrbr
3/JSahhMEcM1trKLUiJ8YnB4Df1gzvBAWKqa4/W5BGV27JEiB6VntTmHUV39YOKGKXSm+ikISjw8
LFDBrWtAhE9jgOYtW0ZAURNIoUWWyuzWc0mFpwpCPQeW66sA+RKd17fC1ltjhowaWSAyQJXEbtG6
I6fmx+bD6q7IdqIEd5YSuWe6eIajW2r2tAqHTuB0S2fPRg+wa8AEXxEun0hfQWdqgPy5Cf/oZqLd
XsSPaoraid2tl0wD48bWkicPXQ4UoR206s5g4VsERd0rDbKSliL1CImq8ukErHh2RLwPfRKc1Dm5
sYMXQs1YUQKM0ZyTBeq1RSQibYCq07pQSrmo8cxR/pJ7cOWRtM2DgrD97IfehR2yrsDAz7KiI0Us
geW8COO1DweZYdt4bsdZ/lBIuTVdmsmO9cMg4q2IOBrH1Bf1L5BeO4bVh53RZ/C52GEQy0gLWcEu
JqY6lunEzFNsridnUF2gA5V1Ad8Pxb3fekAN8UxCNn+kRhEdKeuXcVz78qCJjm4FTmTRbuxJG0cy
JIa8FXnhU46XD6ihe/FokfMBQ1bMU0aX/TzKHL/5gkDarv8YouHjzm57BavHVAAteWIc7REgcfAR
cxbxt9Pt59aafftKU+KpiohXIUTa8a0YxtYWC+KZeeU6EfEwq7k1SfSTyI7H1pd+opwWK+oq6DQp
hRvX838pTYwdc7EzoFeFfKgGvHWIsLDLAaFrH3eZqJkcACYI9kKlUKGE/K+2QaqbAKhJ1F6dPD22
OMHUuHx1dIBTUtqWAmMWFV4HyKYxs4uguN6+pGKxp7YUG74XBkd0btPOCcKeO45jkjb9XOqHtcCG
pbYiZH/EG7RFRuGQOlU1dJX0uvGO31ItW7zRVcGGvRNWhFglo5kzDQUg0wAP4XhC7BBfHlsYXOSm
0gYq587U5yxd1cFJbg7lCWrEn7wXBM9XZ1PbFQKLgauc5vhZsnOCxG6VYMe/Ia09YF5F7Ethi2+i
bwAU7qkdwZ6aEkQ4nufUrzT2admlXmdoaRxCDpyIkiY8gEH4Gf4DQ2qIVrp4VsS3AdxCNSdoAeJ0
BxKCOQAxryo068Sy7bZJ5CtQN0JlrTH7LG/t41VnoemH1FZ+PCU9e5j7+ke/L9j3jwuph2UcI5id
wfUI1+20wW2lAUNha+n8Q+PTwKJ/LXPvl0ho7my42fXjjPLKU1TOJPkcuPTD2Rhbj28dj2R14bJP
AAlmfSmHtXlSmsZEAnIQb4tGQviEI8rJYrKFN8H/MjFa43/XTJMTZKN/tdyrpXTC6nJbNU/7jycQ
4O4x35QjL6ldBQCPOTJodgvCm8jHzucVPErnyR+WMdntRRYhFbD7/lF1paZWcqAkd7wiHD/KxAEm
CLbOHaiC1/HFup5ZEywzN4UMSlvdfKJB1vc4BsL+EoQWbgoOHoUPjYP7K7XBh7P555jNiTviRnpJ
sn1wEli0MG7LnPE2gqz3drNDk7Wb4agCRtiaJELXfgc3jDgufMMbLiBB1heSWCqpXVuZJ8WWoCga
0XAV3FJ+sjFgPSgRY8n4HyWI3XNa8Se6D+MyxT4jrAYIRtcxopl7axQSSjCMo9EXLG8DyqR5XXhb
E5twqOltozr1Bo4iqLLhFCAzFn/uT6gQcZGOolCAaPP2HYqvg2oVQjBtv245qStQRUHXcwXFI2B0
KyoTaoXgfSa0Go8Ufu8MmfOW2+7tpBpB1WeON38Y6i9Aj6ZvE/EL/jHQ0Lo3CvA31k1lxj3/3aE8
+ndkz2uHdMotxKa6cJggDpyT2+nWHuUDoHLMacIoMtNQkUG5J0ZJYpTRG3yovhdjW1qNCWmnHUja
Ji44uDPGTy+vyWl0ZL9NQr4sU62Ge2hmffU0Kj301CBinxZlv3lvo75GbfJBw5YGVcxidzZI0As8
+AHr+VGPM1jSZi47O11TS2Ia/PcUI7w8yvq6e2bnu4yGmpeLR4pJrWSXb6JRm99OvenUTJlSY0Ov
iyhoAleMxIQaQe2x39d18rA52JSJuGdzzjEVgT0bfuM+qlNJq9FGHqlbHi/1Df+TamSFIshlro7A
vOSmgrRP0BB+IfzldnGJ/DZCSOaE8G8vRPRsQm07YOmydUsuYxL6kxxJxfeKOrmqiV8nNaF0XglP
w35vVIzK7kO/FfyPzm4GUCzrWTYKC4cIU7QbU/YW0Ak+RnWixKzsnwT6XHLAO1PjYKvVnRk+VUhg
tlhAB60cF2zKE75G9PsNRGUCGPEfaM5dgxM8ZUMxu3eWnYTVgZj8LFVvem1XUiFDBrqH0jdrvIjn
I3CBDQNECeso4nViKUdYBUAyQHb+wQwPWhxJ6D5lwm3ihe6hb2xkHm1gst02BIbM/iGmQI5QW+P8
RI7u/o/Va+qpQNVJc2sTnG7r+6WqWBYgOm5o9MYHHAc0Gdl8HgHgXhz6x0MCkN77q53H5HVqvkJd
a5qmH9JB8VCworun3xvFHLq8oDdMppKy0MdnRIZZxDHV+zQrkBHZcab2Ihfre7iu5hAgDREbOJJY
r4vMv+B1uZsPqsn/EnopewtQRY7sXw2wO2NECXvrbgu0m6juvMnollUex2+nSXdzEHVs4XNUtyLV
oGNEHKpgU6aMtBhqfcAZllD8tQe2UfXKFjJPUBHokUeKMcNCmKEGvJXbGcrKg+K/Dp2nsTTLC4+L
jQuil4b2ODaJID+5ppmDGFmZSEUyrGmhUcWED7udUnVX1GGsanXNya94yrR1o1FgS/quqzFh7jmE
0H7hRiOIqbap7ia0aIbRt/ALkb6YAuPxzTfF5F9Na2aUislNUlP0Foia7dqcl5J041q0zxfizocr
8EypaclMKdOrWgM7HLmvyKuqxY1r4YmBrQO181/og2ZQ8WvjIKcmZ53p/dgK3MBTLVZN5zQP9ROa
/KKFM69mojoNnRkLmCSkYND0QF3zF1Zsp1U4AjDW+pETrnX26SEa1jwwmxxS3yxhFuEu3QZUBqGO
yqfyPxhKaQjzyRkAd+9ddB30sNdlO5Hp09vDHPzCnmwUzpytStuGaAcifv816VCotsMh7GP2EVdR
8lG39smkFlk76TO8ISytjAFtpqBGfckAU/ViyrXQtaHXHehNfU4o6OQKAh6bB2jmeUIZLNi/xoU0
aymqFvPr+Ln2Pc0HXezRTBq5dP5NdLF4Gvda7umOS9Ph6D1NATtcq1AG/3qe+OU8WJO+JnBSMQlH
oE7D26wQvSGvPrj+MmZ5/QsfkgaNLPWf2ziFxAD5bJ5nczdYuCulk0f6F/1nM10BUbtua2OTHM0T
dZs+Ng8UUSspKQL0nJp7l4ydoDyr3MXVX1mMobmaYMiLsjMAQPSvNKiunEfsjJcACFLCPprFBM7B
fFh942oTqhKoDQltAyi3TapnMtpe/4Xx+GbhULjC09SvWLj3bqyyX6lEmD3SgXp+ET0Yn0/pmTyg
vP+KEIurUn16+kXQQi8NTeE8HqyK6F3phrF0NlQBxrscYSSL9PYBZ0aBXvRY9o6/EZJ9ZAgLWGKI
j8SztNB+WeXgxoDlszH4xJxYbfztRkOOmfYBLB/aonbDCkccWIFvOQJnynnpRE5OcE28/ZHdl5Gn
fFtYWuNGf/AmgNrpw5IFvpYLSvKT/IjfEacKxI3Z1Qy7IFhjy8tAZpeihBcll1jX0HEc3xK4tghl
0U+/5RbosbzmJWczmHT/cAybmxXPIKxLYg+EtBXOoi/0TEDSJjdXOW6aL94JFtO7ykkryPApbew2
UbmmQC7tvKOuN+EPMofTOnCO3SBHx3RWm99/4Oaj28MUqeJhjyhvtE5uT4Qz/U05vUoAcyO8Lt1K
1uKNwc71OIw5xzqYgxDOkRARfxxQ7YETAZ0Ds+FatgDXOJkFtdCqMSFaspu7OpFkx4yF6gRVOige
51ZMRLh01fUfXyafm7b9XRwiD6HzG17dzXX49jZN0epxtpY14yFkkYYTDgZ5MaJb4gfMRHzenT1L
53IcgmIPX6IL1bFnlFRw4cAANNMliC4LXeyOLq32CTuKeB3fxvJzv9xsgFSVQDnYoZ2yD4qNTQBO
BFIb3v2s6dtPY5arsUoEKZKya0RcDeYUi66xwLchbebLcWqRahHqosQZIFfdHlhKYWv9cmF5khYj
Bm8uVsmOxxtVvhAusve/2kFF4iLdBo4yM9K4RcQBCFqcVu6AQeCBHw6p9QQTfChUT7gwLCvzVvnX
7lfEuodkSTa5Jlkd3zsdpt6haqBvDxlRnWF3o3qtAc3eQBRg9b4hiN2GUXQSOwP/t1gQG9yBSjGu
1qZcq9wGla2aPLXtaMn8380pBogD8AevZ1EmaaTCiVjB6fkzonYU1JlLGpiBDmiMKf7Mwkhk0bqv
Ralfq5WtHsHEAOFmewxovtgi22fxeJwPUYeaFYylCHxz8cESzSrUKSoaXiY5WQTi0KUyWswhf933
5I++kaHAudgLrwS83FRnVoO3n+hooGf74iRQLA5S9qZm8skBJwDHDs43lFORUTRPaJbu+sXFdrug
/QKrxTHBrEJHFwDk1EWn+nPKLhLP7/3YokOZb1N1khYQ3ENeSnk6oL/ozmHKjCoXOb0fZvq8oeuW
cgjEbqtWRhpb6cwW5iVoD8moEDA5s98dQFlwnXn4aokXK7ODlNdtkGSAmbu47fU0ci20PH5Iqy5F
dGFnp4yrVxaTxo6JiMfwHle+RyExx245J8BIdOTRn0wAsMZhpAfNzQbZdY66Noguqnv10eI143Xn
O3IYWgWf2DetWZEK4SX3aGKOKeXPMZn5UkMPUC9ccIInirjpCAkk9KbnITmEcgVa/G6/CtSHo296
SHn0QTC9CuCOPjNk0uUVMG1Ar0UpNCm4/j0+2fabf4Kq5ZpHL4DRNCriyC7RzkbR8dHsoQAvAors
cY2xCwxNdhbVO0bHVAySaMh1YJpCqcaa1VXjY9CyEXFahE+gqZMb2gO95+6BaFjoUr65vcs/k68K
Jj6us4wAZU74sPmwA39ULlNk6flqP5OjBE072b94pjcorbe8qWh4mThaysQdPV0LwK0kiEi3YnMg
dCrMbpsjLegfK0RpE8ckXjrO1riZiZV0l5qm2eDEBfuuZQUklYH5U9YegxsLNODwI+XDRxi48fRt
H6ULUu8H0sGUEbu1v20NmcTbGs5P2wUvmqIrXbmsXpWLsTzTvLoUKIPDjpIKf2jBsp01zmqq3EDd
mM38vcoujMA4njFEbC2UgOnwjFDYjaC1PfjZQdFZqTUYEcz1NeyhnbB75hYYi/47lLYYEEiEhk36
e9rNVGAxKk5PG8iVFgLKRp8xJMqw30xNy/2kS8ZUqVFor0lnqVlTCF4GMnr8KUEkUqj6BNH9c4yr
0p+MzsO7TQmAugrZVZwl0BDHEKyjGDa4g3F1QPyYFa/3usaIADgTvJU2mB1hNundLB0IBWow23Yd
G1fG2QGit7X/k2wHRWQYPdm2jV2zQP+dCPrfmTNHYXnwHnrmNZpuHuMjyZdFBeaDYL1tKLjVH/RN
vpi2PglHh9XCriYFCEhah4gOWoeY5G6lm47jDIfykD1ssFCbY7UL+5GkEvfHD/6WADjQ3Q1PZmkV
iiRQUt8cpBwa8vjQ5J3FvaoyPwAx4KLPvFSuQQAENVcOSxFUZZpUOld78mVtyxek9UsuxOPYICXI
YUwcxwulUE/va8CjmRAbrR7paIMn1BBpucD+36sxDdPxVnd0bvxqrSAYHCP5ZPNqxs56Ea++R51Z
auL6bVX6XZecq3QmYVqklBdZ3GSHPtUf3Wt7VSR7P91DLYJtZp5bfANzpGDEbeVFvfmWmHpcqmRm
d3S9nTlpUQ5oNp1XCJLMk6YzKo8pR7Ou88a1JEhEfa/buaKqWL0qf4F6494XN9x/OFpu4BNXf8Ao
Z+IK2Io8rHqnNUDj0Yur7ffDTRDVCveLQhXc7RsmU3qkmE3l4FeX/2FMWGnSfsCNrDjyIFl43VKq
iUkKpkujPbzG5foNxUoOrtYzX5u8ZQ7b6F1N5bS+gSOCtX8vRL3H+55GeC03gTs4jJmIHyZ6Tld0
Pbt6AORbmxTfB+QyokkDGn783rob1j0/CLxIpHHKSmmZz6+/EtVqmXeH3tbvZg90e/XD8+DgZDDV
amY5ZRISr0tOEGByBa/uOtsNKicvK7gi3NlwBC5dSkUSNQ3pGNmekdv57jagfEQ3kIsrfKg5gVsc
Kk/WWTh7SUqeuTuWJYVVizgAN0Yn2hQQUjIWexd3tKGwCvAdHLao8pKBqhG9lscUxftnTz1/3gSE
41sWUOkiJgtUoHXUXPKS9oYe+B54UXj6+oZxXJbxBvdhgEds2N1bh53wfdN4eSFSVjcL5Oj8JYYB
kUxB6Kq6wMT0FYKFe742WAljgVHMDLfraTtNabNyTZCT0Xj30dKF6OqDpQ4qr9szJFZb57X6IhuG
V72KCu6ZsN5ISKs1M7ivygV/zBFu62oF5qcOEmEX5yC4Sdpc9j1bOf0kZ9v0q0oCeV63VGU0xchM
x0hGWBhMe6UbYBSB4mFT15uZaPiEHi8CjhHfQLpY1BdHyj0tN4B8PfxdKqhJ1oB+11leo96f3v9D
disWt/hq+quGrYVrCYzCBV88uK6oW1ObBaGDpqmfKqO6FevcYxO5LfgltgtW6iErpjDoS3noro5J
ycU+zfBUdhiNFl0tzFmsL+USwqv49IyNyxvYejZ/BPbxJuQudp9LtKfFiu2KU3pfcPb1hcJHayj/
bDukRvOj6+ngfQisowRHxjUqMjvZhZuA0dpNMD5d/VKrDH/g9fclPOovat5lX+gedoRaVcTh5pY9
+cHLsVBhi/+1OyHgLPUh9HYkClQviYeMW6om9RYY7yjoGYvaGS7BeP1/VPFLBgnU85D27CtEgdv7
HWq4Wbvc/GzwyifW+KhsXSFkid/ii+Tb1qDvq0sWSCBlkZ0oKZcU8zwGefD8Ex5jjJ10k0PUoN+/
symwrnVWR5kMd3KY3y+qhOZv+KhKHHARcT2OdXdICMLtd4QqITOfPpuvwaVbfBWQGr6ZT7Es4QKC
M2Sb1Le6XgfFpk492TzEbtpp4/BB+WWNhMXIiq7MKOTIx7C9gdt5FWL4IHSCUhTKFpNJnlZAOD8I
PfFv+5kwdF0OQvSBea7kMpe/Aqe++oX0vvVIZxeEKO7EQPZZg72k05FkEf4K4LorT9Syg79AOw9M
2e4hej+ahhfdehxVAxSgjl3ba+Vrp9LEqhYHyxvhlsJh3BYggoZsVRhXJexLXInzc9eSV23uI/xC
yGAynqiBwopqzxlcOLyVM2VXZx2R28bMkqSCyTZ1ilCNSMqpAzm/jwMb4CQvoW8mwBzDSytkVOzj
Z7qv7BtleTqg7niHGHZ0GT0ujNgVG+d4lWizfUgNj6D0TG5uOaFf7rdHazmbaeo6szViS6FdP29z
9R2CMA0BeyD6Nh0EByGi8b19+lgDNXzLqYF40RGnB9/2MZKN1uPQ7lA9LBDyLrRUdPCkfcmU/elJ
8YHTFR84SbdDc8Zqhx0axm/bE3J+R5AWJ18PlbzX1shjDw3wV8PTPhaslEBb5mcRtq6HxnI8OsKD
NUh9LrlVBw4QH0K9rKfJawIGYLqp4oAPXOgnIg+N+9G+nqktTJVV8+goZpC8hAjfAzEmkRtySjLc
c7oVFuGId8qL2E0dw6W7k92IjAOIvjueWXStE4YdRPI6eUkkfL09VG/M88PmaoaeLT1OmGuuvreQ
nSjRcSr2D9W7nXnzDCIexNdkU1LCP24qpl2kwbN+rhziYImanhyBKVV5HwsJMRqYGoEbk4FjWJ22
SvOe4Ab0v8Joil9jU/yG+PtooYOSPvjsXuUpMkBlI0t9JOPxy5GphbNYPNzgXpYetdCEk7ZnKpns
j/9LENcdxjgIuQympB4VTtkjyaoI6SuIU7ki/mAtTibHCxCceXTrrh6J9MU4FtwqSEOLcuVWd+Hg
2QifPbjpeKpadZiPAushrWTwMbwXa0t/y+Fxz0ADSQgWIQMAyFvgBlkMnsJT/8ngPO3fnDqmkVVs
ttXzGz7Z7NfGv3BhgzT+53zOE7afTOoabBDZOt4VWA4mgcRqs2T9JGLlA5w95h+1+PdYOnpvYjM6
GXYnH+xjuXjW9EdC4xssGS2ZnorkNd9nbduXL56Dqyakc/KK6sQ1xCQ19K1J6bjCrijkp8QtRBY0
v6Vy0S6+uwvzjMkcGAkFOOxFFEK51C1ydJeolLIvTup3xeEI+oNdpalmGJZbTphw1WlD8HPGYQPG
weUqcpvO4+rBPwmYpx+nyToNAmXbB3maSE/toh2VgoH+4p3gmQmwa8UlROG0JHrf4t5a46PG3U8u
p2u/MHDYQUd9EEe/YCSvKeuEnmECg6gkiKTu2wI67LfE/QG0OI2KlHh7wUJk8v4vLRHGVeD8EcqI
RArsXMKPhGFB4dl5vZKdui+Z9jreI1jaxQgSJ2MjDl1ibDcqCR+YhGigwsvuh0gpQLDBjdZ8+Cc4
pc0dEHW8aiGfMX0vbQHNgYxYmeTDxIDfwNN87is21J73D++WIYhwHNltTenO3mexQJzMMcRKhvWG
xQXBOKbNFqkzAyC1pTPZQWkPYHJNn8/z0Zbvm0MODdDmiKvzII2636/xEPzwyYo3+ocs4WQQKPVL
Y/cJN3CstkVpcl77VMc4F4QeWoa1Y+/c043YH5kJVg4DBUYknNu0jvm3FY/NLLLfOSa/pvZwVLHP
4EwaT5v6GsM9Icvo6wsx+fwl0aRh4V4ejaUPUwBPd5lrNThAoVSjYya4PAg5RBwPNAsDbSYT0rAB
5rfu3jPG0N70HW2SRBu72CQT3PcmaZHD4l2u01kfOar6cfgXChhdeH8ONo55NmPmT2lNk+/IWeuj
Qx1XnNaLjH0nA6hrXX9H7XmEQqW8SGFl0J70yU9pDeAwqidl+0zDFDxHdtG19UAGy4SFRk6Vlh+g
IneeUMxNUCp83ttMkGgE7J5+lhXh+R3vmsdW3ZUCsxqhYnXE8+yh0iGt9XIHYpR/EnXaSpduVsHj
ugXKIP8EDmBW8Q4O7qiz0mqdXDWQLY2JyUkhiyqtXe3+Nb3VX3WgW7jImsxm49sRADQkmmCDNaVw
t2QFIfdq7An+Ki5Mq5ysuiGzernvMsqg73kbKyV3r2QVI6eOMn9ufeYQ7pUTRNl3hazoZQLhpaCY
Fz9SRT5ofkdaAcQdnFExHWRUeCGTS/yPQj9ydJa3X1Jv+hTznsMVWu2xLkLCCGnWDak7gsgDCefd
RbzS/EgTtyiNkCSwlfPLNjEyvOQbgZOX4B2QnoC9R38BUW9vdTiqAt4iuPORFTChwyV9XU15BcLz
QEKJ5L7pwww8Dl+PG7gk7OOxFU5OGW2ZyslFopBwRZBtl2wrc/+dNa2MnZ1k9E/PovlMSHjxvVMN
92fkofMWXdbGllGCC982zuMX86qu2JqAaIpPHVL0itf8zjJtjoI1p4HbRvvr9Mlcw4c/P0ORm3fr
dJtixOfeTtfKXwIYF9U2r4/+mJubEbBTqlF9l87etOp2YLi4IiEtj1QlKkVX1TPs98ALQMlB0iCP
EAMqmxPkea8HFZWuWfJvRoH/zjlWRx2Dwl93e058TYLMZxmWerzGcUZQ6sSYafZ350/Jz++7ATkL
tUO3KyReRw4xILbWM/fsBZgXCVNj2H9ekKP9LshyWeA0iH//NblgFpxB4HqtC/+yvEtjrXjsrNXe
5YinwBRDDDZ6uQH9fBRuwV+C/eMC0YQQSV8vtvZTEmnVRlvUTl5oUIO24oFCchVevooo0XjL6lgj
pYst5yiQEcDxayX2HoMu3VK3cfoKwfH0cquVLhDcmfNSsFrc6MFnfbTYvly4cpG72x//wqxiqIDs
6rOcBCv/3pzhS6pm0ON2DcdO4TG+AhcHgBLNrInUQgW4Zu2Ja5NTXJ654Y6E/nHrg9b2gcMBWx7W
trV5M9SgQrXL1ysbS2mh40AXMJtiLAmzVdUw8R36o9Ssz6FBiozWRAAPmxLvnRjJm/RxuV4chymE
CaT36NxHCGgHX4JsLqj8AXSo/J5W42DyPkrDi77jb7lYlSqRoOI2dfLm4BQAIHy7+8rbEOoXdQly
hqsJTR0q9zKlPIwcO8ryNob1ivBnB+JfWGc1RsAZNDWA+Obt5hIu5gVi8EpE0U869mqF6b5wKizF
NjGGLgAjHfCGKHWbxkKoGHwHat1jcfMjI4mkSJzQs0ZhJJPUUP1xYi1U4qfDpLbe2XAF8uVjs2LE
cJ7Vcwko8zRrQPDzmWeQXE19pl9gKD1niTumPCRrGPq9ZzDuicFR4uuxOhUl2rOGQIH9lljjOQGk
gNDCZX9M3WVMklA2A2U/J92qQSBJcNCwQBPvlDwapSK/opdu1Rq8KYSkrKrUqmLjCUg90oXyb6w6
LTLqzOEiQ0ixBpc+tMY63zoYwC4TP21BhecYoWu9lpdEiYHqmquLyDkgRizJan/lCIwlwqtQ/ij+
Xl11V5T2M28h+eGqaWrXwnUnI7RhO53CMxzN6QyEfTrHQXbkARYzsisidGhsEWhZOk5CBHKbDeCj
gJ0sb4SnceSHShmdO+Ch5gd+OKliW+K1f4spiImqLKWNzaP7XXhjz53e4C5jc0khxw37sWFGIMMK
HIF9ECcEdhRSHftqv5OGtThjy4zNYDqVHSLy6+BnkLrHSlWoBAT4lUucHL87Y6yhDPoVIVpICTSM
MPvjakHfZ7iJEES4MSQRMuoyT9FgH2qzMTC4g6wENru3z54hXSJVO4WKWn/QGv8Z7riWExGj2GOu
b7QpCIW7LCqW6p/+PAcUrqxvLF7UIA97DVsk4SvcITZ/1y2aENy/phwISQBIDN8NHx8sHouJaj4/
EZLUGFPhapAyWf3nRWWPaEe0CibNYBKL8wHLyRHOjQUatMpRruIIM9i+EYj/zsAU98IdHNorbgZd
fsZCyW0F7e5OGNBj7t9Sk8cim7amB2sKA90lcLntAz/lRimtEf40H1HZLDCArj9raC5PUMi0jthx
GQAN0RsCaW1l3oFWobkSgNi6W5zQZEA3tRpEuOM7EpA0sMl6qZD7V55MUTqkdaDjKkF7KS9UXonK
4mNWQyg+Rmj502M0Rnd9knjZ3JkjnR8ZK64X7ODNRTaJS+d/qhfw5g2F+WBETOvRk245ZQmw54K0
LH0ZprHc5nKrdvXxDsDJ2NuoMKreih7+EUln4Xt4NcHhVPmP+/w5RnxoiH1Pw9U3P9/UtOgPANwx
kQXaP4xAjqeM2KjApELq/aV6c/nlLxK+1KGehpaCMIz54vjpc/LhTod92wSQeVHhGXCXXC3X826V
HQcDuNNaRd9w0GejrlqMg7kuTrauT2M9MY3TCyUhoRYcpvhCs06/rutvW3Zdkg4qJ5Z87kv+KSPY
4OEx5fVAqbr7Q2+zG4iPiYpYTc5fSWcolQe6RDDmYc3iZJ1BknKDvTKpt8L/SHY1ZaJ6cnQJeHcW
9ngDgZ949LcRGWM3+DzrwaGwc8mki3qu19Hxy1kgU98GfBG9sn6uOFZfYYcm8lyl9awZn4XlQU1J
g5UdWR2wC3nriCXoqf2c2lOCTg+fmZOp5fF6KA7uVnE5ug0TG3IB6SixqV8MtkyHLPvEee9V88rZ
a7cFU0L1ErOzWjDdbm3giMopxZAmayqJXXQubfVqqN9wGT6Gm5QxjqV6D0D/FBump+Z4D1zOAlZn
RyMbxRchO0/OKp2li9aouPpseKrzJUYeAecEVMQTKtV506XLWfFLKAj/TTfJV+PIlk9MN/FF37xX
VJTWApMGIYqd7CrrGosuSsPwAat0MziTgDj3d2/FnedHmOHtNQNRgvjybLLYz241Uw9jpvncf7Jx
U7DNaBd/OwnvnOopTnkxXItTjvR6TO7rEglwCmTWbWpOgB2xCsjC3CLdMAQpIqtUAFgp7BdOpqeF
xcesJMsjOc49kTj3CWiy2ztmd2TVFnGFaI0KpUfqukSIG3pwvike0mxDkKIApwgz1l/+eJIVIYWn
zPRwtyHuZBMTTCuazbIg2gPjgJC5IVLufjZpFv4b0umx41ghiHGf4Zs2M4L9ZS1+GvH1A2VqmiWe
EBef8uu32kgaSrMcxLgCJ+k0H9zzVphen2S6GtqMn7GxrhcehHge0rF3DTgeAJ2PeBBBbwJIJY5Q
MVl96cfeRrCV6FDCVx+6hPjlAoyinXJ2Pp7UOKXR5vlR1Uhvqpfn6LMflJtOBACOnjYTpepiYexV
8oSC5e9+Fp6HjrCasjvzDzM/HaE9M5JkbYYmV/YymrHTVXHYkcPOFq+i3bEX2j3uoge/2JFCQVNW
dURDxTjWOH7kjHdJU8EXz00shynQc3ANDy/cUhro+qDGVXj2F+McY/2FUm/zh8TERm6E5wmlNdWp
kZm/IxcSszaycQy8WAO+IDVPcpNFys/r4OKw1XdTpAOQ8VMRQKWsTWjqBBwcbheQGvM69q7A9SG3
aloJPuRK+vHKdMieCDhhoKuAUu30WF/BwocSdQfHhRJjwiQGiYDYTF/FbLgjrwclFlvC99Tm59Hd
alXsZl9TBxo2f/c15l/wn/X0Pv34p7NC029iOwccAkuU47vTdC7aLn5nxHZSfeGtyFGwnFx5kJ0X
eYgH+7E7jrBJbsvBOPfv6mNU/2Irn4Qd+uABggKR3eWUmniiKZdqUY3ZBy7OHmr9ecaz/u11HP0Y
v/iEnyNGBvtngg4LLOQeMrgJKqkvOsStA0Bz7ixf//i/HVu/zoH5/dTOxQJaXjHcZZ6L6N9I+ZSg
adqK+aP6Oj93RtmheSxbVxqsAGka1QjEpF0oi61DKPFLLlYFeHggzDAOKBcAcQkNofab3tLKG56w
C+8fB0DXKxJhujFt4wlGXYpb7Cj3UNGLKnu3iel/G8KiTgcHNVNXYQRyguKNzPHgpxv+NmbnItMk
YBW3KltlpmcNrflOhrA2N6aBu9tehWq6kI/3LJkeYZV9mZeTtgCGfL0SdDKTApJ5n8vw4VlGIbuq
uVsRfso6aqK9h1P4VxSN+ueFDKvi4h9JppDv9w/BjKHB3LLIHQHgPRRLePRjG0NWKvVJ5b+2+cqG
z+TbvI9wV6xHFEZSHcWcQTF9QyTU1qGSVNVejEElZ4hOOx7JCIJ0aShhu2s2D6qNu0+6TTgDYyXX
PJ/TW2/oVSf7drpkLI2HMMn3l2NLkM1L5jYydh5Lli4rPVKiod/KgieC4bteSs25puprjLAt9ewz
+Sw2r0VfkYNfaSzHTmDU8x4x8/dBl3HLiMsbFMhwG+Q1JaHHvVNBSZZsd7Yjs6cMyLgUoOq4H6hR
O2Ger4VpyOIaPUgy1WPQbecszqtSZ96/iLY5o6JFvdqz4cLzmv9BvNYponBONRR15wixLKkRGlCH
V7Bunp/cmViXA4dqdmrayeNLnq2gZ/6+Udaaeo9V/VQVPbO/dSI0uwhmvloV0OTthe455DCDONxG
8gNyLHKQWNJSQnrccCbcnAsJhhcuZc6hQoZAhaZBBp8ZsfE7ku5HiJNXvhrgAfRjuT7dqQWm69Mz
5FKwNbiElnr4I/F2ceK8371GAPaMfqkSCmobJDGNrAW8qTlMD9x/ARPu0xUnCXG5BDBt+K0DSJwb
8MOcCbGW25LyaADhEGgfamjNQOuQ3UD/qELnCfW3veeSvY2jdEbagA7pR611m3fkCqwsvc0rLkL5
dJobQOOkCA0r0aAT6aPRe4yMEyc0PG6PrjClyKgdIOQMcocDSvrgCaM3HI2wbd+ZHrm4zgVWvRco
8+FLg9txMEbyxA3DTReCNjv8tsp3AlBzcww35Z16/H4Ff5QgGhQTTAEsdPyVUeK+7mTMS1Qfndx1
Ubq2XHbn0mPadW9/0aCMj4YiRGNEMJOZvNBzdHBOtusVMfNZo0/0rlH7ZLX/87RhPFDR65xoJONC
/4UUGXxuXNI7t9pUPP76fk1E1JfUH4Awb82nqxJ2bx8yHB9EXyWnnj0cwDP3iRSR7XmlrO/EwNL/
WiSxPmcBCVGTgdG/FMkZGR+YBPQorSOaJ6Iin+3YMxqGOFR8jQ1tuTJNpAllKS37uxsgQGBvJ1bW
Vh44rx7mv2rOacbYEdzEmLW6T/gqBuZ0dbZexZ8GirJxzHg0r2eUpXCZBtj6MZRFwSzremDuG2S9
JPgmTGWC44w0vc++TupXABcO8I7YkPOUcwiavWLpXQgJPnZin2X119zuiqlUeNonpq0zxt5uQO/B
aKDeotKWmBiK3jJRP5gbbrmjtPJnjEU+m2X8qket/bf/0ExPAK7/BPjJ2d9ZJGFEbsZ6dxNhJR58
ZEgXtwdM/dS+VhKfXq5NmMFh1E/JvfjpCBiUieD23CpkXci+5xi+8P69rdlkG8aj/4KzW70liYER
DgbXYMhceBuY/GbR28T0p5azyjv4OOrCyBxE5GTqj9NPDlNbtX5NU4FOVxqbYlRHWJZ8OJ8G2Tt0
5gj55k8czUpmCDuFoqlJ7ZsyQIKQNEQ0gCGeAhNI7As5KGWigl4I1IEGSGQ0NSmoT6JL94eyhr6W
KLPxBbLJLptA5ZKZY9x61aZKB+jtBBplCx5uamTdSQ4y4bJxjqo65wXrMkLXUOam3yDdm9902DE5
IREHYQyiNCPyLpY8CU4Ktx87gmr0s8SVJvkJedxHK3FLgh+Q4/VOPA8sd1hOX6I9YrV83BItqUPE
clqbe47uNf03t5Ub7g+q4vwp4mPzBNBmjl//jD3CYE4hzKuwfy3bYrUD6KYUjOMwE9RlFMID7BD6
5RkvxEzDj3/333E4JWhXZYRo4dX6FO6+TaCcG2OktUyDCl4RJnTXYSpAOqU/8y6kumJi1vcDUK7u
q3kB2fXEnFF75gRIFuuTMGykHjzaofCktFuuNuoO9QXW8qaaF5RgdBvLlixzcEEBr2HNANchniUc
blkMiAmsU/oNpxfARcvuSQwHjSYjm3svBGkyoVHhwNy1IfCV8Ue7qDDGKNXjvhcb29/QSKQ/A8jP
PEGrlO/X0ezL6qFttbPAInw5NtOL5luCHcNnbWjVweZgCImJ+PRkSQCE+1RlVdTC0f9UjJuhsahH
kYsp4AU88ScMsAF7Wn8QyHpk2CLpdTiyK5UJubBF2nTe29JPvtYEFH1JItCp2W3oNuYuabJ+nEak
jf0c1nT2Y/BdC5C5GXo875FU245rk5uZcH48wBnR/Hit4KexpXgGMfQilEoktU9fbmOSxWPDC37R
UK5RXKCsMN/SxXMXKw0RS0TCpJrtx2NqtC4Xwf61z8vEntC7ORoIe2J5l2+z6pZmeuJ/ysR42fuG
rE5GqgT4skeWzg+LxBJjSi6ABwuyAJLbEpzh8wCRPLIyWhBbK3yRYMEgLd4GbGMQ+uOlIoASsfnV
xqSR8beP6Bzqjj2R7QM4CpUp7khbdlLH5+GpAErk3Z9jcDSZlNACYvyy0WMIXO+9312R/CXhIxSF
+9oHpSWRTgg+u+w6zbTDi13omL4NH9vFO9MSZkU7BL46dPYOf9DSXA8TB8WZMBh/PGL2eps9PAAA
zItIBoCoOU3g4NedsEeZjmMWhVROL6nSNvrFfxfRgJYRXu1/cYtyMg+F2PQhu45+LfP4/0V6pNDM
DSKbW5szEKiulPN4ja4n4SM/4fHVG4S62vrnAMETFNbZflPv687D+A1yrAyclkX1cSji5qlhWikI
a8tKjYpwNHP5Ipym+JCBpHVbhh84hcKzuIRxenQlxGLiE8EaWYst1SzpXeunaef2emnnllYqO2MX
l28YycS2VrGKyNTJEFe06/6+mLRuIIyBwZzdTIB4VP+1cNmfdzW4x7jKTI6kLgV8C5479PEU0wkz
ICX+6oKj6JMCo4Aal56JdcXANWYhlOpvx8LjXRkbCUzBTZtJyWrtFw9ZmLpaxkPKy4FuBJwdjeNY
7uE8LHC062E/PARhI3qcpBRqFi73178yw8bMFU+BnESyk5DOIJEGPLDMWFbPX+Djq/BlB49zdwBw
8I/0x9XOX3wJz+8xT2oKKfnkYm8bYeuRWilqxA1iqJDDqNwAxa0tluT+ycUBMwzMNYwsquIT0w8v
/IZsd3tLE5u7+Ain/zBkVo669X+gMoYVHEhUNNWOV1xSwJHaagaY2TDED1q3SDYkBO1D1Gq3IRSz
9pjb4eK6LAkXBet/SaMmb50dY9Re3gqTONDdbBnVSudL8yjj8MZ751JcbmUpcNia1ucap0A9H9Qh
XFXLGocvBWiQiUidzWz4oWUg0ubWoRGlIEvn7WoyuhTwVkQkSy1FWTLgCRohLsmzLaTg/RDbPEeU
3l56xSBG5WSDQJfsJ0QyvWxOHE3nGMBOiqvXu4heHDyI5umtRWx5T/iz30eB/3v0ZaaBhFqp9pRQ
uCn3AmAp1GDv6Wgcgr36lB3rn0DnUwrZCWWokwMWo7WLugCX4GvEkai+3W1977BrGBmJlsNSdCMs
2yNJzNGE4D6Z+I5N1GqjrHeLeyUuVR/ujBEY+fJuNcd8gVymF6JzrB5ff7RPFBtpi2iWysNGVCdc
Euu6JldQqyaV2IPW3kLLoUpYLnSycpl9h1+9AOce0Hflwhbvx7tuIuuu/1kO+JEpRvL8SLmy/blg
N0XlgAw4nS37n+2CJcbvh5i/3tz/rg/4sJZcrTABf0KFXmmU9QG6XjrRs5HoqCwva/J4lvRR6jNn
MfIFZ1ztnp3EAKdjANbmNjzJqehB814yuqjjxxU3CX01kbaDmH4g20Y9wriNHsSI1yOkuml3+i6B
4/7CnjhDQQ8S8UbWKd71lIYVDRx/pLPV5xJkPmZjH82P+ZiQwlMIVmFLhP61olHN3vflCb460fdt
hF33p6kMeYmCGh3d13u9hcIHwVXQm2q6TfQko8rm0udC4n0jXLfPStlRKdFXPL909FX8vOo9Tp+W
0i5lopYNHEbHO+FJ9FaI7SbRFHQEteNJGT//JwtH6Ykdp+QXQCkYedriBmTrUrGs+LgYrujaj7Wn
7jyCwtQb8Vujgq8ZsFLDZ/Qol8FtHxpHIQMnifjJ7bIJxYl6W3cQiUuaqrVC2LAgFIgk09ra3P9O
M6UxAiY+NJOWCkRN/UDVM1jkq7rN1F30Hnd7Kg8xMoH5nImNohb4SmRxpzyZTZhHNxe4LgQcUDh1
KcicEsCxvSDK1l0IgO/+qR9+JbWBmaG+sN7orq5m4BZn28GqEW0+lbyLcTgcLjjPRJZWfje/4d0n
edGUc/rKUngLzbNI5ktqeRT2gWyti5N1nMBhHR0czFTP2JlgfPBVagVR2rVulxrVc1s/F3M+r19q
jmJYY0Vgl2bzLsCd4Wwyer0neHrhRE31URjF4FCNovVWr/orTgxUpori0EbC6jzLkkdp9NBT1Fpp
XW/PH2gxGzk1No2hJ03pkd/DAP48HKlzwb5BeJKpQRQQ7aCAkaOAtt79bSY6KOaFC5wG6x8KKUjS
6xNSd2pj/k/nU3WR5FXeAk23eFurJEn+TkorqPaxcSsdoZVDh+xud0bVSHCOPiHLKi1MaT2N6MNa
h/9FaFffapwsfgqBV+Y8hHdEw7uSdUEjaMZGr57tolgBVK8l3Sx0vq8ZklpZ/mabi5q0e1RgZE26
ENcI5gEnblVRWh75w0gPyup1tJQoP2HVs7FrQcgBkfo6N0t974PGmA139VVYQwfwdFNvMNEirlCC
N8mQz/71EhPXdv5FnV0BWIkrxafpx1AGckbm2rh9cetLdUyGDdcUboKxnp0dgMctz+kIViCdFmgI
vZsoPNnmGm0RkuRtpifUWfyvotPJPc5ryVXzfDaJmXJ7pT28tvUJD+CGhHd0txhS0acA65Gonj6F
fk/9m74sTATLWNv5OTPoazm4u5vEio/CfxcglFodvReitFeJ+40VwSgjzP/OtYgrYtylmpzcvGBG
xRN+ZTJh5BNfskyOt5gni8Pf6Kv/P0XisxesTReJssxnjwUi2Zxx0EQHJh3Fay/AF52lADFV/SQT
kCePW3sBm5zbZinIdUpgJ/h/nxs5VUDlRpxL3YJXPZ6Szf9bhOgnahVdQk7Q73L75vpOE2LiH18h
vVGIeKyj9rHnDMnRinN4DNKMyVbYG0BxDYj/0WnMS07evq2HxFHYETDyZLX/yaPWfe9fVffzFxm5
dfiiu9qE/tovPkuZvxOWpI4CX+UR+CL6/hB7X0moeDOXmVKUkSFRYE79JXxfeVm7RDpDCTWX4ofR
FBD+ot0IcWjwVn3QqRvdctVTqmJ3835Hhho5KjdjVXeqRsi5LRcUkkmUfMEpB870mNvHgdVgVBu+
3uGrnBfHa/AfgZ1mFaxErywiuS0RE2c91FpSxKGaVTM8JNW4ugGJtPoj+i7+8NUedO8Ys2yEb1Ir
IxAHQ4QwVzeVsJObNlpbpXQisfTFU6TsJuY6Bghgc2sopLa+QP6zMb005yakQrkjZGslT/NAUyGQ
KRLRI7eXZeo4fuNgv8Sw4aBJ77qZUGoIaEHB2Ix6vYLrdPWecyR+O3IpA/2543futZQe+xMVREi4
1HiaVHMiF8VsRLN69ikuJ5crxIUYa63MhishsRrvdvfkx3C0NbPMkUsv8fIWAz9SP7s33YQevx/i
Te6L9jMOGWKpaxx31d41YlXbctp8P6i0ic8029YmtMP7C2hVemDvS6KZ0sA3bFxk79oT6Kj1IcB/
SmZefhTJeYwoFwCIaHPOtbf4k1Zn/tcUc1oQl1+lyC6+FX2+DUFN0rIzm0GWbE0UnRuzHqsjDWDa
WSUXSreYZglXPtGS31HPaxmCSWbh+SM5KuYNzkGZfcsjNFDliIwR5LDWX7vJxS3wk0rIHnCEs0zP
VFXSiGDOzIxSWvNq4AYVgKQKv9W/eyS2LUf3ssR8Z+LFbNm27tdnXVRV8WkHOnADi3D+XgYgugN+
8csCa494tWeHc7prBsRkGx8X0O382aUjszQLMX7aenU995Ibzv98ZIL29MJ/GAUdq6A97mkDep7N
9KUNigQKpGlm5jfr47rVjYp3kf4NvMwSlOr2fQt2mfwupLIyyod8p00roz9aTfEsSwtvIaj+SoJc
pIu4EQ8giC4OjcuIN3n06i3+eiaMGTl3OkXAJQYW4dzLeTecaM5y901aMHGACxVS6rH5ew5ASIQg
gtsgwBuOaH17j0kO0T484b5UpRmjUzuW5EK9WBzvXWOfO2lwC5ybUqVuTgApdwDlFaViyT4sx+tS
WlVztFzRvNDf1x+oxoM/LCJQAa4o4zDe3EUhXNI7IFDAwEfEeToczvxIQbHBB9kB3gjpYZ1dQERT
DFTemspjTqlg1BEIffSbIa1XxaO/vqKwiIwBLyne3pNtwS22H9iENsTWPwGQ1e+e2VcecaJZGE4X
uaEepqA9k9ysDYlVq7gOuO1oGhc+yQayTFUay/G9Y95p7izrcDsQ5KKhLwC+tWZjBiJrLg5UJORC
dZcjIbRIpCfa3BlzhCR9Y6JpdrUzUAYg17VlOk7/KVaKnJAGUohDCoVxuuKeMnWaJntldNCGXOic
hRCp6FNn2UihXZcKZauFYE9jdendzyrGCjZ7hYhNP1t7LiVT7GJR81RA5GqpJ9eJ6YLHvTsjH4Hq
XRFws8bT0vpTWvRVuHsNu9Ho/M+XmfVWfdUJAxeiHlcTT/KM2LLSMp/t9DiZod2pKAMso1kE61rT
tPZFpAdxqjfVzUXSry2F1N2RGP1MHF8IN90K1a6khmOz86emxs9r7vKzYA0AhECoHjlVSsSXe6IH
NnzVcNzcEP4Mc8UZKIz4/1zVsCBZ2k8/wdU/L6wWZo0GTP7srT2/Mvoq1CGr6KW8v2yH5DrDvl1j
eM7jRqW+AiHNLF12xz4iCZl0Xko2f/zquGiDXPsV2q5deGZ3Xaqb9sGUj0MsG1RePJMReV3HFERM
Eqy+PD7jklZn26ZpVG3qGjuoo65wHX1Y4TCKx/rCq3F1rcyV+q+T6t8Y+3p2q4m7F9oLZUHD+QFq
2BgRY2+bCTo0/MItdq4zHa622cAsnaOz4AxGJUiPGJfnChOso3Ul8B/61wVEEm0ckoEsKy1sOppH
9mJ3YBQPUa2PFDkOwvaInMZyJiRLMdzdU8dtUMJGXGVSPmIQFS9qePrMeiQHYWIwwzCkFwpRrSmj
NOxqaxy1k9qkyhrJAmS3Ghki6XpBEgCHDGNipRNmJUA8DKzIXzAFeeMQ1kn9CbXenzngt7G4GwtF
Df/PcmFwe/lVSrr8gZG6GMCOv+H6e8R//QmQYE3CKXqcFH9/yPJKAxLlFFThe5w9jH7fUbK6lPpT
nauBXH5c0VfmGBINd2zEYEmHdQK6H7VPbhkdsOQAUj8j9KnqpXBD/pI4fbXYQaJCoLdFgYLUWllO
m9wv2cyyA4Zk6yMzN+v2BcuE9zh6X9BYIP0RHS+BErJ8Ly6t0AbMfg2jljJPSjTo6B91+BFfkj4Z
NRU99MmW4uAkX8ySp9Zd3tpVBSp/x7KgerJN9UJHPZA92eGO5Ezb1CuU209Ib4LxWEFCtvnn6rOp
rYdZM3r6LxfLR1D+xQD2tyeV5tdocpiDw1nyh6f6ZyKKmcaGNCDR4LGLBdQcHw8/xo+6JnnvPdwX
SDrk8SAZRkAdCQhBSbdt22uQUgbnDv437xTO/glK0JWK1LOYc7R1/u7BKetXicJyqzPeL5TPq1Rk
CHyD2L3/3axwQxRFH56QGfHF+aiGSTA2IFKPRm6G3UaQt71Jszf6V6s0CoS5nilIn9HfwhDZT3CU
uAFm8y6seSTtVRrazjPwKLqIyOJVHwOmFNNu/BSq2UGgUE0TseSNvO+ZSXXrZDTaRjGglmtkCFiF
b2S0631DIojGytCC7HPKNGmmAb4JRNnbTn97O9kGZohHGH5ZFMKHZuQwwdFtyL6vqXdqmSf6T0JD
w+US6Q1HND3Ect1BbnVHYmbT1ZSv/ITTRV85il7PKVlNvmSU+NtmnvIrkk4XkWoL5u1QyGFFokwP
ODSRgImwNH6eH4PlbvE52PcYEvvj+uDTFWgV5yhZ1HbkfFduSLKgIRuMlAS0GJLBUBilNNJUFmiC
za3twyHW19UKodZ2SrK1wGIq/z5nd7n4fWRc8ZvK6Vftsf5HQhaMo2bbkayJgxsXg7X6pW/llb3l
ZjYSl9h7MBXx5BNmWzVjJRdHrDZap6bPIrhi94E5VJwTcmfzA0I7uGHPXMe9n90FxxpD4IRADGMh
dIEUkEjxt/gKHAsPtleqwzmnHng/DKSwrY+gEfrhDmtqO8rERftj7TthqtMUGhIpeMRVxo+CYvOG
SKHT6saLvPAVlmEn8K4QhhHM4+ASQwdXnshws4EnwJOV9fOxI7krxiZSlmCch45SHLHRkwWfryui
dghoEpTYcQzAXkMZJrO6nyxVFRt3CKFvaphOZAF93OKLrHUoSGMkbNFC4B3P54C9iAl+1Sw/TCCz
qp68m81eunL/feFmW67XT+AJWqLam98l8/nzEIHm4FVymgYZGuRnLiYawBVyUjShwwyLKAV40dAP
ux3Qw464I2IRgylF4QrgQ22tj5FjOLDiwtws710vWwkNzDbD4T4CPHpnE+qqF/C+OYoUmuS0Mfed
19xpx+sdBNJ2TkMyiAN6sAsjnTeMMfb+LMBhSm43NTU0fjLx3wnVZW+b6AyJwODew3dbaSt9zfr3
I9tVQV/p4UNFiqEQpxnCTe1ZpuW3XwIl/ECNCLa+nWkJQ2BR2aEHX65tIagFA6vUpOc8J9IF/PGW
WryzErSDH0n9HG+2hEBHPCCKQBQIJ+zQCrrugeCHqQs6Ui2kZnl20U1JTWCbc1B9u8w2G3YMJ0e9
0+i/q+dm8ZM/eTEYUmhe+SabEKZEpPWa+N9JAqSiTE/155VJ03gD1WBbcvDpIJBa2bYu3W6Y49+p
v3rOTqMq0+yuypykSt+lPDSN0fpaW2h++B4M9wecXEwz2NiHXNU0/qlasPZAx2H3HO2tBoxuVweF
KP6hnNfSdrl09b+jazSaR11b7qhHRRBrTwyxxSwXZi95vyCNWzHGyUyGfVM6aGOZ1rttjS0crRpk
lVesSzRdsz6qdhPdNsuRO/OyH5NEQm+Y1A/xAnXhf633y6nF8q6blxENylVnRSADeqBN0gDreyo3
vu3jQPmIylKLTP/tJRJe5SviJjyZuxYULrC9TCju/U/0qfghabfUe38yB+V4FThmZq1z6C9SgwbF
Hg4mt9LVrUwYglPlrQbR12OpTIGOaash1DEZQ2Cvx+QaRYzCTKSPB3bjUMLqXEkUjDJIGq4/GhTa
J/jdKcvtvma7Z7hsXl/APyN7waYzyF9ZDhnjwrZ/+gvC94fnHhuSAVe2Rf1wwpGWI/M4PKZKKCq8
hljjTAOoULduHJrhUbspcEkB50Zgm/7KNmoVMeTP9Fk7qS9im8u73KE2m6rcbO/6eL4SrN5J6L2l
9nl8scntidVyVJb/Fu4BqTVasJaTtRgj3Gx7/HgzWtgJlndbQ5IBMB2P7iHStbIkr3ppGBYx7JcB
6tS+24m2wzRbgODqV3M1zQI7VW0WfvzwaVhj1EtE4d7QhtEMw902DkXtB8ittdRqcq5Hvoekx8hc
oGRilaV8d7C4qkACRgfnFDXSDpPlsV37PyrhRzX1juN+V8tjc8/nYJULjLBKlDa2UTrS4RZKZePH
SShusKzYeb6fFL1/6m6nlBHE6bVs9mNkGXyYOcgCyONRUf3ZKDMqE3ISK6Ug9N7lB4uJt8nktfE/
XArqc8qLRCAqijh9GSmrzJkfwnRJNpQW7GrqXAmirQmKusgCfsRq/6o8CV/Hf1zkTSlXUYi7TRKm
H1nPiU9ukrgwp9FDrTYKW8ZJdRhPgHpVfMkM6DVUeGzg/p9+anL6hY/J/LE4oQqZYh1DD+GFG3Y6
27NUg8VIPnznMUTQcfbjpRg9kEmK1QbGJQFklLjxfX2P1quJ23cz/9jJHvayDiv5c5sK11fbJWw6
nZa4qqPn8KLUbS6nI5NTWxUWO0Wkis9A+QHZqvhNTcbFyLQDMP4B1SY3bnjgIzgs5nDTwFr91L2C
g50L4DZ0x7i8ia5XN5Gbm9ZxdArjHcGHzxcpqGyi6AXmXf0xarBEaDKyfnXlZVb2ldcFUz3GhAaG
ssLa5JO2qPFtCgPnAe+no00BMLFoJvN+/YxpKd4CUABjZKATqNxSqUkwKORDetZ/9fGokzv5gesW
VYrBIQpZBpL9CF0zhIQWN9zFFM/AkXNn/ItR8a1dskNUhdkJVX38hbbn9JJy/QGaIOE5HaIzCLia
jwLqMFUDCvNLWsPmINwt0n7JR4J6MCPXaibt7JZVKobtXc6HhzBwTMiXGMF9WV9vtPBMIRtBZ+F5
p191egv82LiJOvpYw+zg/Mi/k2FmKZ+54Wlewd+OQUHLJt2lWcPoDEEOVKTV3PUlMAJ76/Fu2pVp
AZGGI/gafLzUU+iC1hhlkjVa5el5m+4Ji7yZW/4z549B7uBdcuy/6HltNHWBqOAnhi8LFiFg0cZd
Jxvmo6lxP9ZUEBjynqhUSYaSAFjL4/bsbb1QOJS6q9070ehjFoBGJekh+G2c/jy7AUm3475a6b1s
fZwKroiAvBAnZRPskjTLgYIWlQNjewlErn7qyYjbgKfO09TIK1trDbso4gmuYqGRk10Dr+In4gRw
KxnnKutnWGMzpeGWejbeLubEZPF1311gqhbT7DmnkqwncGWhchs/SBUAoRHQL4RE21ESOW9KMuYY
5FYV1y+g9CHHDEVgQ1UqOgwPxWHmbHZy10OUUf7tdC5KVt5gf4zuG9hkTv39H2EKSZUWNkFuakwD
t4BNW0/p93kJNFVTjvKnUMU1tIg6pfau7Ki+mP2WrZb3kL1masUsF003R4VGbkuEKxL9idRn/QyC
VXBdNv+GWLFVWEJn+sH2Ds5XxAE2TjUBA9aEE535wgfsi2342TYofShgXzOUiPIO0RxfhmofRX2z
+SB0FtPVB2oGMmIbjsfvaB8NHsz82lwJuO1WDCmadNlXOyRKkV0a/+MUx+pJemi6H3ZiJlOCy3+4
tsOcC8ayvG7Fx0ZiMwT+IrUfl/7OJYcNXMZmwhf0TayFJQK4pSEsNCxFm4VfaakArDwH3/VvFNzI
S1SnedES4BJuuvGa5Q+6K2q0WJHNgJiAkOER/4Fk8NexBJa++5w9/lvn0fG7Hv7/m+gLN1XxIc31
XxSO8v1pid23G2rt5pN6XkCAfym6miPF27tQaMeILN7G1w/GH8p0jNQFoerBGjNlcW828wH3R4zD
6HhPxFF4tOUF99wadi3m4LywLy0XAQblvbTjMSNzMW1CvEUj3Ky+aMvOiwRmCRbxQfj6XoL+6yBl
Q/ZWbXNiGskwuZB1vt5DxhQIhzLj2052tL/mWPAKAOyKPwzNYxeMpFutAx+6G2Cj3DnmvPvIt1Yr
Dcg0OHn4cOM7I6kPf03cVcPGLueSIl4GH8QbPxECOG1drVxrilctfSuq75OAuTrJtgOkIa3zPi5n
N9ZL8BzkeP8efj3c8eIJRi34NgzHChr6DDRp8FXuJpcCt5TbHQ8MUfIQy1kWnvg5XbH8zA2FpQRS
9NNPeG3ysJpIR1cuGvYm8pj+ZA2AE6L9me5qg18jIi6cDlfOTE3BaMiAaNWNWh9Zi/g+M5+gpaOm
G3PUZI2GPGPJkDWiUW2/4jcKSphsBvNUDrNL10GYsbH0ZGJGKv+PbWCsRz9ldrFYtblfxMtBrfvH
xXp/lG4v+JbduHVRkBzlpgJ/jQMGcY68GkrgGVmEZuIu9yrChhwU4T4lkScznsGGWFIUNufxjdr0
miHqrmS3UFZPjek7JSIgtlhBj8z3hlsAOk+2nd5ExjRCxqmFcHtQUzNFsKYjiPct5ZwrhRvuntlq
tiIurwWz37M97rC01Tt+Bz6TZlAWnnymVtFGxeAmPcnRtayMMh6bUEg6cYiyvCG0T5ZnNtIUcUkW
kcIAZN6LPYY3aRNW5+BsYuBcQmVyUEmz5KeOQwEUGBVB0UyQ9GkOGUNgwxNfFqcE7qWg53PDQscm
dsMesGREM4e30xf6dDxTEa17sNNidyZhG1LvHjbyY8pEasPXqwEKPjArot3UFFnTADUC4lznfDQV
/CMwKlnNUjfCmfKilypcJNhyRE2wACP8kGoJjlLa4M/0dwzjWCdp37jA3KORy16oU2Aeb91mxF0O
HkKq1MYFwKbENish7blMU6J2J2PQ0mrr9HBNpntJQ+3/pxktd1G20BwoJdeJZGgDdGUGXiCsUGt2
gMJSPpmq1FS4r+wRh/hdRQll/2QGkYEdSCue/agvNCKOCdYwQGRdfpqaHjCcnJzo4uf0XWXm08P2
XlvJlRAX7pzrYujISy6VG6R43/Vv1JBUC815XrxQqSyqy8hm4jq60tlUwXPuKWXNpt1StzNfEnjU
nQV+0kfgnN3LNWjjOgWJjmpsFXTpCzSxYa60Bu5TpNH9Fvve1PqMOV6mTblbrqbUkv2eDsHBRf/p
9t3cd9VcoNDk86qxZagWjoNY4iCdzBVp34pXVaFHcekCATUX7pnv6LB5GtxNNc0nCbO8s/LaIVgh
x1dTLh0rpm/2bzuq1WcmPpQUfPkBLdK985R6FAulAFLpHty5jjfKK9FoIbuWProZp9tAbJaQT9r2
kOPPalhxh3Ov76XAgY4Dy8h+7Lzi1f+IwrzF9fgArGMl1DpLeu/UFgIeEAp8HD30igs6CcbnirxT
hurQua8s3M9GjZZlRd/UDLo9y3RmtEKz0ghCK9jvfmbGq4F6OIs3Zsjl77XX5wBENTPH1voyQVFs
4SvlivhJibjQ0viTtWAD6SIHhKrjjpVIS5J5Omf9VjRQtrXsX5ndcK+Kb5xVjuB2hrCDkPnbiq15
wgzZQSlE4UFpjF8itH1jqbQ8pThkoZtuUzvyZWrAgc9m7Bq8LcWdWnFSJmb8bAp2rj1YR1ky+CHu
B+xA6xlUS4L97PDeJXtHUYtowIWsmP0qfocELXWWvvc7p3wcUYF1gUGyW0t9dGv0TmCMurepy3DM
Ih098IPYJIXnaR249Hi+ATO15DcXLV8P1/oGX0AVN9yhRi8tXE3Akm/k+M95q2hHdl/zAKsN20b5
JJQ242LEGYg45jzPIsA3yBCaoxPadC4UBydw/EYYU7ng6fGA1b7/rLGcjy9w4H4NauPHJAI3+/MR
ae7EytGErugpHsUcE/y8lWbHPVvTr9Yafl5h7l7p5Kge9VCbJ9YdOi1gHYliYF0nEjSnhZlhODge
Fb9/DJjP8rxWfLBzeWDUOcsfJogvw+7MIYoape8cdq3FT48WdnhTAl+dCd1gfFOcVzW1WRYXOQpL
PkFmHmdc19bg0mAaBW5QqI1nE8k+D8pyRRK35BchNiniUBNomeWh0Ezkugd7iYGENEO9hx7xwatf
P+/ep/YG9OUWdu0wJ45Ko1aGYCMMvHzm3ftIwvKn3YNQoQZWgsPhlmutfBcGu2Gj//asQ+TFR3BN
BaA8rgzQxtAzHGgd5os4DCMLz9V9y39krpXcOXjoQ9nMDZLn+NmaIfPUJ5urZmjMLohkBuRu9mMI
xa+1Ydl1pP2BvwaWH+vPAV9sa3i0krNCDUGv7xQL6k+wsjIqkuYhkhRRE1nyyxlcecUsuXSBN99L
uqvqiT/XiVOj+tyxwQH6zStZF/Z6kK/6tlbTygtOJ72M+lIa3G1jB0HJsNI7sjQR2vpfqQ/AEfnf
tmerQ1Vf7NhZXkfSfFSn3+6F/HaLR0oF+N981IuRswi/LS8wYl7ksFTZnnUm38tW4/MUGnvWka8J
yEfEGDm42ptGYliBP3maeOXqHBTzO1mX/Eqsl9d2MRxQRN/D5ERklns9WJ6DfAYcRWH1xpV6Zebs
CAbozKIjoskoWE9N6uvhPI808/y1Ldbi51AwzQqHVNYDxhRdtmHYMflphcr1ZETCfQZM1/U5/oEE
HDaxpBOCqJ7LfI9f5gv1Y01DlqebwNaUfRVARjMtkyojKk9esEt4+Au5rGIrFTqWRswU+U6T2AcP
2d2kuRob88KKO07e4I4bGAp5QngPAjBoFR5VVAKxi0VW9DOnlxMkdY4dIbQ0KdXBLWaF0Nkn39Gb
Yg5p0v8Gxlx9yXWpckrCAKX3DndLXxkZwUb7KG+H4cD7XrisFSx22i5Dc10Dw/gdA17diHXx9WDT
UQTkqD/JvBl+2q9aIxxyW8RokYpv/FfZQn5HsMrmCgiJYuGTBDviPqJPRdKUIZwxqWVdwNiSbGCA
hg6pQfHakadsy37A4klPQ491BoXoPJHhdSTf621deJ9qfztQr3Go3a4zLVIxTZ8eeNBVeL2Lkdd6
M/BFBUYthoiN+Pt48xpmt8PQbSHvyo4Ua5IZNjA8Hn/qSB4BSui4kwdGA15GoOU+RIy1WxhYgp0I
mUXym/QNL77T0YtihRpl7jGZAy/z/souXYuhqOF1nNUDkWNlWPLNUJ2/5E4xcMgl530LciHx8jR+
lEaevZfV8lejGUbRnqmd3k60771TSf4IH3uLqRqZr4nqkie/g3N0KS4crMhwdD6cohayE5Y6sF02
Rjdc8SDPxjp8Mg/DdBwoM35Da/M0KfDX/MaTspSdJuXxLMFpKNNN0hV4zXz5wZhaHj9Zx5UzCzYZ
CjQ3Lji9Nf1NloHtjDzgBK6fYY+OMZQUfNuzXQ2JLupUSen4r56OjJfvcg/XHcQxLS84I2Q/3G/x
sYXiAdpTZWvQxpeDTKHIzo1TmLQLvPxvZMMzpR77abPF39zCWghverAq87GUgQUxDYtl8Sir0bU/
P8eEjJLH3G4rZ/TjlDOdgLPZ5oJkKMiRrl6DvrR0UC6INGg+IjiaXlnz2d8Dmv//Y/qd4bsFn0bu
GHPyCcCAyoFkBfGEYw+s88feS1LDUixTQRU9zuMIfJIl3dC+XMhusaNlRDcFN/VtENLzRDYM3cze
ovuSCzIC17wZSCUs+fTJmNz6HeQ09UX4VpFbBS5cZxP3MfAWEaXC/Y/RdVpT5JusCtTz9Q+Gv6RD
cVHo9CGgJ4G2+Bnmdmkyzun3FsugVF8uKakgQ3WVJXr8mxFBvmsrweL2rmMegVEpqvAw/CYeRM1Z
Xb6GJc8fex44uX/o/KTAx+WtzcixaWjxvsUrravyGj11xfJl/4KCR+OFU9sryMfFOKh/cunsCZg5
5GPxsW0g/YPlN2whHJsJjg/O7qeJfXi+4AOGl8dvHIQ1fEGrE00zwPsaPsqcqouOjcdgFpdfcThe
YJJGyH4QHIMNXQ/VAD4IWZo7vmRUDyT5BVqOmiBbkMXPk8kI46anqdMoZE4q5f0JR2WDFCu/RNbU
62k6O0S8eMZcUa3km4ltU8lHb9zIXIXzBgUBJaSntJHV84RJ0/ZF/mIXdUgLDlNkrOzoGu52AvOs
1FoL2GTTJDwez7awbwVf/A5OYszuB01cO1PF8Rrkt2xFhDQo/Zc51Tt7ShZ785kCl55575KliazN
s3EF/Ad+aNEcJR84m4hOYUZNNCWzvIhzrMpkOg1ycnKBpLu6Tq07F6a1DIT66BcRPQ+YaRFiWQgo
06BUeKoUA4XYNRMJTEGEifKTaPgEYFeT03x60943s4G6iqMNzWGYnJ2aSNvqtPGA+osbGTCGauWM
M1SEgYvbsAPVHAcVtgq6MrbVi6eHGeqmbaVVgsWAUGn6TgzibvHbmgbJynFce17735ezKz+0/dP3
vdiOO09go/uVl4RdGx+Jkp8SxFjqCgDz1VuQ4+3zp484uW37vOuwzD64CA89LMov1WaU4bjqviXZ
LV5rlmtWVDc895Mt0SD0uV/0leqeAwfYa6nVxY+S2rlxDYfA3UAfRcS3vzQmMab+EA02y1HDZXfR
jT3Nnci2ikaAdbDMMsavzt7WN8qM8umfIC73hmJjFGcuPCBTMkwaAKQydarly0PiY6QDOHelberW
Bw+Shcob3RE2rwAcbf0ewvArYGGnuJ3bGLqn6TYy/613pipjQhWk8cGx5StRKDklnmTgVn3+6GTD
XDd+T12Vvq6CNww7FpYirHTJIynAicaYemSdRNlnfaM0hggSgk96nYKX8tFDxmXeQOJ4dsn2S+IS
8eFfT4xJp/iTZYdV478JLJx6mpZQGyAAi/htSrnVqJeLMwca/+DVY40OtB1VZeCSvFRRyE0oKQFQ
6R2+fxk7U0UdH6Ux+yLJuODgNAvJl2qNlGBuoThwIg4FPATODBULD4bYSZnsGrb08Yi6pc0yIguU
FhWxpoOwadCRZelA4pS0UbVeOeXntuf7aLhvxyli5RGcoJoasvEDJkQJICIDO/kecEYktnpLKsVw
beTwpd2BceUoMU4uUBZSmJ904c6qoSzdgu1MAcu0agNiO1g70TmxIVDuLNTzutK97iwogzXvZK+Q
G9dkduzUU7CxgBbFV+7/UyyWCikLRvt1vmoihmq/ivRfC4ZiD3VHk3yNE/n08nAf65Zyb5bSjIEL
dlvvXUK1ZpjKaZn+71P0QzAAwhnuB/bv6sCEN9DnIISlgFOLb8POGKZaXAXu0Dm+j0+V9TmF09Gp
oG9qPXIVGZ7F/wxM8RadDUvTCQ7qze0cnq8MxzE8M8FhxgD7p29iVA5dK72tBOWDWH4VxlcvUXxn
4tQJlQ4QwL2gOZRRU/TE+yqwin9OzhykHvDimfXK1rmpgcVMP3ulpwe/ppzf9XA0qouuGx86+O9J
HsQiaTN6tvNi5bx5gnLWph+i+KdntoIBn+OJdaJJ9ZQLPfm6ZFh0sG3pcjckmL6EyFSa20EY2VHS
p1HG+WkIHMoxl1PnzChNz6A2IVtYSF9HmI6MJpmIc+M+6XqgwaonJA3/RfUd+4kQpLxxsMcqtWxm
XpCbEmSHt/xPhbBXde1H+V0k/vEhzpsAD8zmi/BH6p+wI9hMiiJDjl6/pF6WIFkeYgEeaGr1NOhR
dMVW/ElEXQreCdodOghbPYE7EnIhRoczZt2G8IUNVn4jqiNg7fB9EMZRsSRuMl6jrraKnWF2WZbJ
PTMYOQ7TJcpRhP1Oa3IVkIQSpOQpGs0PlHQ5XKrxLN+zl87VBxV/prPNnF01WrmtLBW13Athevbm
WXJdfeBbrJvjnnTA9/9k+k8LhjAuyOdJ7lfLpakRA/1lroaMBA3GYaKs/Fet82DK88/8quAXmlR3
+j391QW6b6giNvzplzARPm2rPFF6NeLc0iCSQOu999iJnl2JXlPsvoECFiXQ9UU0nt94IWmEBwBm
AJVYTB5slFWnpTWrjcRDy8PA4eRnNsJsWEPRcWAD+l2EeBDpHB8JXYNcB6CVRKYKD7C9hDu55jng
Td7gih/AetoJHCxN7xOvEFO0ZlGm9sHrdBLXy5p5SGiunVZGydfOd44aBAnBooJTYXmgVe3TZ+W6
vRl6kIxE+XjRJ8CP9clDFZ8RuTMSnB7+K9EJ7B6psNrK1cDMofJRg75f9Pk3ZQ5HZ1GGkBhmG0HX
CVoE0maD0YiWcTD7UBaDb+meJJCANmRBmJ2/7NMnvpXXmTnXY8NucgBbZnB/iY/UUBnstJiyD7I6
1tsb62W1CIKMXRuVWzMeCS1F5vPQ6+1MmnSlwjAwtPRQNgO2jUYaIBxpwHVvWsu58EmXeSruYKAF
IKHDz6zYKmoRG4lBLvb+dqE1P1ou/5SCVkZsdgGWmcXV/kMC5eVoszwQaTVVexjNFqYQadkGG7eZ
dBDvyicqAF5jS2GZxS40B3BB7aANSxGpGdvaQs69g8d0aj8VIj40j3yTOTMD6O9R5TklZaPWrP9X
N3z/RgaUeLx+J93XnjGz15eKrIdr/QGdMJkegNVAnK0rWnhMKpgAfhFbZ8WE4/kA5/bYweIJ4L2o
klN66TYb6qE9rzp+12yGF4BEckEaj3EfT3y4pVQPm13rZNxU2qOJqfrTf8BG6d4C5TxhvoLc9cbX
NMWOJ8TnOLsLy2AYIAhZoAzxBQF/rNoFmnrAoze85yV8htwt5iWW5QNf4lwVn3mOUn4ZoNPr9h9K
KePGIgmf55Ekj4H2ajD7KFT+xYgsDfurwviwBNisdquL6eSZT6Zm5J9RPA37Wv9jJ3QKp/VIvdRY
dRLLCCPGg2BIMNEds4QWy/gz59WRkn2Otmf0UG/jfG049Ztu24vJf1vT77MVuIUSvfd0Dp1AEH6q
cj59CcDNwG5SE1+nE6roBWusogtR1n/VxQNAHvV+i3mCyn5jSfsK90M63wcJ6m3x24X8eoc22j8A
Wn97w5FmJZ7aN81omFn6JF9Kwd9mhnBSgZXodxtT2ZOL3deFM/F7wa203/d+MKQTHnivMSHZQ0sq
uLMZ17+OhpQmWTu+xrnLIerzo5yr7V/LRUL26g6vVbJR7eTgn8zdrqQdnkuixSHMb3JaBQIVbE6a
TZ04HchUnbvhmh6wOaOaldN1ETmrcXLNts9dILeWG4+zbxEKpXvz9YmjHyT/+lKYMc/pQ/8qegtP
maPHMAOCUWhQOmhViVV2O9UtkqKnc/VpleaiiRbs8gOPXK8xFlfALxXl4EQQ7d4D75nQEs/O6ESe
goptijSahO9/FP4yswsKaFl8za0qucIHLvObNttFucXY0YefymtZkqH+A+LSNo2DqsJOpjgV413s
YnRoP7iN17k6b8Wg4MWyx70aa+KVi1489vuNE0fbVU/NGOwXhJHwcl+edNHMDUAO1CyuRCnFwRqX
lvozSTY5NcUK7KfptXz4TUttgbJuLVnc3ReM6wBk2uggMOuX2ul1haFAF0kNVilLnkcSwJCUsyo/
5X54X4go8eubJCMdbUzQGGXInlig3pcErx2QHHfmeCbzxa1FJ8s810FJQRm2q4LS5BGiTbgrYU0q
lN1WIcYFh7NjED1luS1Y5uFeIn5K1tEp1xcKVZF87nzQBwbXnPTQgxj5s+16b3QsUeDC0GnKWx1Y
EBIGiqyW218WaKPxzms5FcG8D7JP74j64PqCrTqFQci4yVG0hixIQpNlOHaBKRAOrnVN4fmy3L71
ZDaueZ0uJ0fyN9aDHclxThj2j2f5ej9yhMYAB4R7is7KsLalCbG+vSGsqLrvuqIeO637jTNBfo3d
tXOUUQh91LkDWgK07+l5G3Y3nt4m0Z3cbFu9J+4grHnbqx1cnKvNjd8sFxYWwt5j+8mZRrBEDx0t
bpF7MCUHmKpPsiVRYMSnkfuye2onoIiZWaoCMb/uDxTA2vKag4y4lVMWQ8XD8LJFi3w6B3USwWE8
YJj2p+q6mu47hjar5lq+HOepwDoqaQ1eR4ddqwqyX49RUnF5JJSrSXvDdlUlxDMu7uiMbEupPO6q
bIbQgSk5LXm17VTeXGveUXUPGABq7iwtgG/JmZOpLBSWspsbXjHcHIzkSEoCsSTm5vQ0XLDWAcW5
jlx1+AZeqnlfIIgM8d8u0HU0+HV/Ks39BzE5bmc98YH2LtOYzUS01YDkwe0NuxtHerxar1TLUueU
NEaz4n7uSUhpNp7neviiW5HzKw7fKcddPIT1+LBxEtWk99W/bZBYOUkauK/hPuo2+zSvKQO7it56
Gxe58l0CGjHmOxs7I6vF1iXui7jFM7YIuH+TQG4L5Fj4mFIoU+GcY3Pi++M09VrLKBSKwiuQYeoh
hXLKBe0PQnoZDe81A75PpUeLr4fZfbal7Go1+tMLc4bj1Pl1dJsnVjocAizDcO33uBC9WoMa8gIX
nDKyw324nkUQ6FgOV2jrR8Wm3u49QwrifNhfZwr7aGwQ3/xMbBTkU9hnnG+bli/gVLVIr4PsNKu5
ZUArOpqW/REDizpG7VQ1tbVaMe9U+7Gfcel8wxnJctt3GJywCoczE5Qf9PRvuePQqPZfZ19I/xDc
kEM0B6JXfQFf8dIgAHfcPU8ON/kaEu2APbMSk8/+I9GtYMuaRkTicWUGGXam8y4h8/8XAin6yW/i
ZPIYJhGus9k2oUVSmpa8H8qnVqg8gRmcpkECqAjlA6z6IVNfScfapfh16pKDghFv2jKGiP8AjaF3
auGes5vFieFh9nbn5TFtorXOcniNJ0Xyxm8sEEB7byRCMuIYP58O+Je69e6m3ymuL4SbNKsLX0c4
GStIp/1zyoXUmVtM1SX1w0VZVQ7cuqJWfxLq1OG9G68iqTRY3Iv9gqgAP+/cjfp7upeBUm3EHJJR
I03HtrlmLpO889+XCxiGcSNBkpXsE5HipXodrRePlf71bvx++73V9A19hO9hARFXDYXbUPwTrLwR
2ztWoEIXOHrD7+xJOKdw3cQaQMBMMxi3oTCh99TMkUIZ0Ny2CExUXirLl0WdGWiV5m08g+rvVvQn
Y6KS+Tl4oEF69mx3NzMVx2HJxQqjO40TXupjQP95E6OOpypbUJQ5516RJhDILOU+qQKAlAX2jpwk
8+HEgSkynS+a0WFBIXcW1jIIi08G4Wb19s7YOhLbDkb9xDTcrwoLyJ92MUN4J2OaN/nWw3U1q6Yy
tis/ek9WiKT0FaCY+KYSobYFqXYq7RSaWajeHnD/kvHdlhe7Z7JC90kEwMuCqLT/12BbVQ92vkhV
CcNmM5YwSpmUBFnrIdWx9RMLnLaU2B241q9UeTOkCMUROmmJ2YZcXUh0+MxTPeCtVK0E0IDVuOsf
5XG5hDPH9KN4ETG5NW4rQ9HOOFAzM1Q3L2ziQRw4CsY+aM6uECy08c2y23mz5SO/wNy8ZelYsAyW
4L6qhcuNsK1gWChjJXd5dPQWWwJqHdE7LG5UxnX29RCh/BI7oBnzbVrgASJduZN7UkR7/6nZPnn9
XsaWv3uD+I1OOF82IRCSY0ljVLKNGIOTOh8+ZC2L169lXinLOoVrY1Ok7Gaj2Lmt6w7+59MxyubN
62tN6CCP9sshsZohsF2lrB+5BjIssInERQ3V8attdUh+nAnLgpGz9Do6QRx9S1U0kbUPHfvtAkQc
I30pWjK6ujmOsgcehiQV2c14pftWLE3lJeKW1tNXmbCffj42majyQpLE59vAvpM36Ykdbm/13tbN
7APlCZqEGHK21tdumAOuX0Rmqh7j7eBWoT77z1nYIPtOH4IgOhZdRePf0//5Gnc/HY/hL+6HGR1c
6G9iovRHmIxv8bi0KEd8JC8F2Ij3R8/Ft5r7Muw8bsOUzjVNOYs9u273Xl5xKRYhw2rlipe2KTk6
3btOVraHn/Igp4cwx8/lewbv+V3jp58nnxM+GgQhfWujRj10n/b/l1Qn55FbhDw/aM75jxj6rGcz
f+Y8gWGrCt8rov3O0KKrO6+MDA37qpob2zm33mHFg8EUtHQONR9XfOxoE/dkNeGHCiGsy1WwW/Cf
xmZJvgIVeZw5oCnABdrQt4PRmcE2vhTFq4uYVbXpMKx86dBr4Fc2/iWnClbGNdE+G6jXa9zZGwYW
EGbq1Sf29bz7GL18ZrFsMqA3Fm5wTlas1sTBSI+d63ay4l8C3WjZIBjyoCSXeSK27Z921N029gdV
kGmSk60GJ8jBuuXTPJPiImZ9mZtDDgqrH8spd1cG64OQjJWIlFIgpCmMnFygwepk9nmFGMkpN2So
l6s+ml5ii1apZ1sPNAmuo5RJx9pjvQyibZ8qCK/kxDf7mhvspTQWt13klqIFUr+7xam36YG//uqp
QVn44eFnqcBnrqutHhb0OhuMOdGD6k7s1QDlixgQpCEosfeluETBbX0RGKsvLfMQVKSfSpvYNuDB
wwLCjH4bpwMegchlp8/C1ls/1w2I1VRQf/7qav0G9y1yNr94+NK3N01MDC0t6d0qIMWfBOzkfoMb
5cTJWGbZE4rLdTiqSJhpHu3lxgWWATkb8ESQJorJDGr69BGsI0UxJv+Lkh0z1hf09kWaoYBBc9lp
HRUEXuN4fiXorFvK4jdK2LEIxyWhbySZVtB/WgMiadrsXaLoVkjYPXaPLuYB5TYcmFy1mxwlS/Hk
x80umvqTYO/Jxv8l/o5NaUKo5DAoIV+P0F3XL05hc9HbQHASPfEfNfB3osH9xTEsZR2xwmAzJdMN
HJBox+1dw60UzLhyDnrb3BK4rmGRt2VkyFYCOQVrFgAwimUVnM/fPgNPFDrbsU4ndqoNN3ePYzGk
8FX//UZX+PTP2pMSVyhdVvZRDejFsHjreYnY67OyDOW921ubeaIEPc09Q2ZGrzlgUud5iWPci2kP
v5YMkMhVQxtRu4F9KdFT/QMLC3tX0TxurHld5T6z5pUXJS9iy1jPDoTyDBGTzuluSLSl2ywYuEdV
d8EtwF5e3GEILkMehWf+F5gXdft/4o1g1ut6n1dUficD9rQ9XpTjQIicKGHDf8ckwVJIaJRPJefp
ztmmwrfvsaLvd0avXHI1K7KXYJ5odDlzIxU=
`protect end_protected
