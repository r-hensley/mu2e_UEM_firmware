`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KQLJVYVmGDiflEsZv4ToPtNEXcpB9Qk1VrCLnQrMLQjD0fecE8umcR41BwsmHX/IgzXu9LeslwJ8
acZYsX5KZg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gc9DWuLlGRPmPi/qwrCmAQk4l08nPp5uq0LmjXDpwIHTO+UknlM3NCJ3BXO/eZ9zhvMVhUBSOP8d
5FR8138ovfR/lrbFzcp5MJEGdZiatPU5psnVRJd3UztVAi2BLrEwPoWT+GAm0toeJ4SZ6vC9tnrY
bmXv8z1YYf4f6xIfLxY=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NoybFKywXZMCNVUi0sw/BUVWrBJtld7vcJj4yV2SPBjFlpLP9sclOeXgsu0KJDDMzDbNhGSFLvqW
FhJ+tnG4NUYeoxTibpxJo8zal7tuNDnF6c5a3loQe7mIV8nm5vz0dmAPphji4n/EE4P1yJtfLyWC
zBTaXHGMHn07JUgjixA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eL9ZJ1BKQdL8n+R6/6Wj/NaLMJ6m6xliLXWdCsGgDxmw0Lbp9ZYosyTg6pUwcCIqvG7zg23Z2dmX
4dcxzk6IsszNtd2NUTtZ/1nJntaqj8TkxpxDLTDMjNCVNFEv1Rkeja+eXvZsHjl3f4mcytxaqthK
uWZCe/Uv+SHGu+nssXjkgSrrRxgkx4FFneaMJki0ghXnVkBdQARcksoeBLfOhh+IdDF7Bx+Zosb+
+HnsiBvVwACLbDB6VB+6q4tchk6yHBEUCnY5haYTQIZHoXyDURQ0xpoN1DqaoEhCKY9PmUahtC2n
BnDBuRfnQdZgyZ7gG3vnu/l8C1fxVMQqglld2A==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KdWDaG0/KEl35DtOIuwURmpLLCw4h0iRaD8yrFvLAAeRo35+FYmwMP/Fd3FQfVYbnsOnr9xep5kF
r8mbKU45oYIwd5rgJP8s0mXxdT46PyKF/0noORz0heWm0j6jrC32lGnK9vcl1JUo8W2gzH63SlG2
Gh6wW93MuGPhIO8iNUHGrlYJLMZe1vAFwWQk5j2Crah3/JvRdFL07bUA2D6W5Rhly/q1MHEArx2k
wA8ioUuJf5Y/epLMt+jgbzpVsQ3eN0YceM3RuAy98/64qSjD02CKLOT+48fZPwuONrJzhM/sXxFG
C47SLWRcyu44TDPhYYScik6xwgE3qWrF/pbfbA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u8SFxk49AKyytSA4GkMRlrqxWhrrSpJsh1+9VlyzLLcpGGxm6LDafc3Te45IfZsDDNrsL3cCTT9w
OBLlDVQvLK6nk3ADxk3gEHf7DCFnnsI8vsGSer/CPlg8jCRPDFNGFj08kCCkLfCG9weEflg6EEY7
FL1g6VhfIoapQSk6sE9ZLNmrUJpzCdAR8JhIQwXmuXIanq9UtAWJM0hH+rYTW/hTMRpscfEqTlg3
6vj16nwf+blIgrPPshGTpBev9l8+YN3XROCB2iQJPveBqPQnEIViW8KJljardr8yrud9uwAa30Ru
AIA2ux7ireVcI+NW1Bg7fP1yRL166coWDoayZw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 765264)
`protect data_block
F5o62xFcs2VsOimlRv+tag3JGrDoPqDfLEpwadK+BLDJNVzTgO48xgpWRexFGIFmYB2Em/GGrpc1
Gxlze0o0zdDy0UJbiIOjsXiwz3Py1XaFlwduhUzX0+uZpkV2ivBr0Ou/7nOMM53Tv7jirRe+3dwU
HgI3OUpCWMKTipxBwF0IqI9PPzRtVVelrAnqQDGU/Usyd4c9e4Nn+Yv1izEdTdtCCvyq1Ik1Pj6Z
Kl7PgSqm6bAmIhmiXrb/jlHH2+Y1FMpdwG3Z0l5jez7qNp9hkk+clrl4P3qlpIWhVX0L+Bt2i+7L
EzOo56oQga3LW7odRvPs5xvslanSfy6MT4fKyERHex85kZR1c77OzVhRJ7pFu5+Kp5OCL/HMu62h
iXirIovuEPrkLw5HRCihnOIqa4l+OGC/Mzy2PbJDgFWQzO5ROsXMoE9t3yH2vuylayCLDG6ubo2o
P//6Jri3geXsX/68pXkYsipAsINhUqr5LtXfdXY49DqjM9htn9kxHE+tE5npBccGRhTUeEyMCvGi
N1WDNRDVZ4G/EnlJJ8SaZ45OF7JzHCgQsWlJ2zIeyVzA4qUbf1bfhknQiH4oQY9oiygFhbVE7s0/
3Be17YVJ5CWnbbL7OXdy5nrOeDvDn3Y29RX8VY2xOkxtbM2Tr4djVKjfgQ3dl4nQ6dWYKoSrvHo9
WEXIOW4s+hQp85jrj1IOFDNSx41b3ZvzsC/B1RRVMahWRmKxkwynl50ly8Mi81LsJNHb17JWmP9r
BbukkMaEm6qHyOgJs7XllvYeZhPNpHalLCo5axvlEck6g1r57rPAMVHBOcQXMuDDEg/yIzld8BvJ
TPMHu0fY92U5b+oXjSRRD/oEzBEy7vv7QhefyfIc7JOj2guLATHwVgSZuxocPu5G0XvSZ0VBM18j
niI5YA3IerTOyrMV3PxeJeCAqvYwl8O9PHCH0neg6vo4Xodt/wjzsLZXvONEgjWi973TzH1QZnJ+
GaIvz7jhp23OyUBuZht1OTW4A6ymxI0uwTJdkaQfOJhVZ04ADGpKmivKqLStXcQQO2BBMODPeb1C
J8xlkH9rVRjP8UFouhooBMCy1VkzRmHqk2nonjMjENOScfwF49IdYPAXxg/wk1CWZl60lfhiGLy0
lPOUMqtxW8uBZiEYxQovSX15jxClSIQuPXECt0/V+quX0gtXKsfoR5zdd1oakDT+n6UZWIxFhCMf
zZaxd2Uk6h5gDL4SvnT4O+eL5wxobBvbOo3DfLhBF44KFbQCf/2eWy+xkM2QeaBWcAIS06Ny1b2F
K0puSQt4k3NYqSB0H3cpdm1eZdjGFzbqPgsbGhZEZB3iIWxnpbD+0yKK+Vm7LABD7R9lyGAGuk2a
D3E2EjBkGEZTW4oD3uxvQF7X/iGNFF/KcnslVBUvJGyrhgpR/EFOmR87Od6g3kwWOT0Q5cYW4Len
1Mq7U3bKLjIxK2CPnXaGdQrahh93CIzV8GHexOG/MFH//eGgxj3xHWcDB3fVdCdLu1LQwGooHsUl
Z23cDB/M1uDF2gDMrggYEZzjz43b4/k179oBeI/zrJMzl2WH+Ktw96N7ETDOGbsKzuh39q3z1PXd
iUfz5f6irmM0YPkL8Gl25fxQrVm7wKekAfeBk1nipWRQGIsG+neK+J7sOXfZvvkwfLCtP6LJAKx9
cjeuNlnk2U/ts1hxmGaBjAIAdT562hrwN3a6U1+E2uCq5PIpSJnVaB66JMDWj0JMouLVY21oeaZl
zLpor5gZ14huG5N9vcNqldY0sSz/WdywmKtGuHlgmffheLqdmdlhYuONTRycqeR94V1HLsTD3uOD
sxV6JfEoV8QUSOsXbu+upfN7ze79zeTks/MamG9/BCbo10Aj7HOKes3E3fDPz7JUDKvdZLXFsqeZ
t3G8rzBHuwJ6Vh0ckaWGr80TpgNBjW/BJgyDeJ/csl24EcSPk5xYxDmjVrwvYaiA1Fgn9doiJM2G
NkVLv4LZF2QzXbYHIi7TId1EMExWjrWLNBwi9/F2P4x+I2Ltnaf5dYy13ksrmFtE+rLxCGK7OyjG
xpnuCEjasawgN5vWnjZE0gBhlh1sC0iSFXWktlbvK6bLK3GsMjVcJFZ8h7SRuRj5FU8Ihej8kMtT
rN5+TOGqlfoagMyeAzUBH2+Q+8V0oQ8KRPDn2F3IbCirg8QTvHdJct4lxk3vh+iLWTXNRP8zQSBt
Wh8j2TBfIisXags6VRgUNwaw1632svqqYb40TRcYUg5PbZ9dVvasgykBLAoabXSUo1qiOX0zHBxS
518bl2t2JKEu9mBMdvEj1zvEx87SWFuedfDApF3v9ihvUUFBvI3rSFqJMTfSEAan+FYb8aDfJYPM
c4kooTlIYYOdvGZVMHdv542OS0V3d7JJs9yyBX4XUILyDMkI2vhaB5+chibpqKt2CNPqTmh49ehK
IcutGAVcfFraRlef7qBrupLrFWU3IGoCCIkBzitoHhmha+qoAzzw3Z8DZL096hoSRIy3r6yGHFEj
IcBGO6802dz9QHAlw4OlRIc5g/e90q8gY/k7A72nexBpnnELhqv/wLYOrH8O3pwXcSwfTtg+bto4
xSHJxfwAPNKTFwcO/gqUfCQBfYTlIENDqF7pF07t4tHByQtfb5sZXF3UFNIHuzE6FGwaDz/qUq9E
/usp3E5ohCzwyoFBVMS/eqPU1j2Xbdqle76rOulsjc5qpLQXkf7Io3t2XqU+ICJYCmCgNcT4t0EV
xjmMirJgtHox2Ug72wGcGK2EiujV/aBsmwlg0P70cShcG9/JW1b3OSXtoAqYX61O+ruVb84FA91O
VhFRO/TLPJ7akGnZxRlh7MVbD+z4KeAZpySAKi+K5VKzS+3bDd1gzgZKQStYQfCs5rcVNPghumQf
LsL3hFcfpOwqAhuJQ1YOV17L7cT/FP+4389dPlakcqxjxM1nzI5FUATQcg+Qnn+CNjfIAN/iTqyq
zXNK3owNG793ikTGW4JOuS/ew7ROlxRN7vHKlJAU4VcAtQT8q0KBx3UiPtn31FF+nnO/2pCqxg1H
y5etepqHkX7Z6SJFShdsH8HNHY/U5eLGymN4HLgaAO8w0LaSTzEpfx82DvkQRm1HcDNGbWc7aoeE
eEL+79TT911ouwkxJkcRAPhI2pT03kg5ch0J1cmIELXwE508HMP5ljwl+/bzUbo/WhWVuVlk/+r/
RyG+xpcvpMM73/53nqz2shtWlGWM+WaY3znNWcc9VW0mRWzUDSYjQlnRVGrRm6T4QvCoKfDJZ/MV
lMdxfWFQGmyP6uNpt0SwlUIKVCfyY750ZEGcoyyeqMcusKgjHUFYlQT6ynEbiLIvSgcp8UQQAZdV
M0YX0PlboJE+OcwSK1JIvEtzt94C9kZd/lWIXhNia0L25IhMOel5LQoPqZ+zDa5X7ounKg2DBaVe
+/fQf5+DitbTV1ndBViTozNcZFqeWDJI1RZxDQQUJiZZHuAqm/0zwVCuduOlXvU3hSn1tIzvhYk4
TPMc+egKpDkzrR1lvtSRbV5rV7Jse7Mg2S3aLMijEOwO//N3kEKm76bNKBv9pX6BPzwKa8ur6vPY
qFY9cB9n9B4p3gX7h+xpUmuEqoQLRYoZjUv4jgspKD1h2j2H1He+vJDZAlVilA/Ve9MW4k/r6HOc
kyT6ABjrfCHbu0F5ycewwn6AJTcLoKAWTaRCVeWaRNiSQq9VJLlt9ga9AFFgA047aZIbvBMEBBcx
5pDgUfBV7EVA0Pc6YHcekCbAWWbxb9UomnsrdLUV50ptDiSe+jqXVgdDwdxhVTZ5oChvrIOxr0u1
Hw19AvHIc+Vq+fXNAp3hLC67+c1m2yGnlu9vxruDBCN8f8ympaW+ISJXrLZ1RgACK/AsQpEo7Sae
MJmMaAMKDAF4sXe+DW4aIt2QvRIbYPPhSYnqgxvzWIPDOYzvoQZQQWmYaA3cVrSLWI9iEq75CHlo
WuI3eFy+s2ufLgP/Ln33xO8jCpxRBGAmr8DuuRyj167Nf4zAvRuCHplXb3JOHc40gPgZDrL2Xfzo
uzIOegzw+cUIxuFIilfqtutX3uwekNUxVr90U6cawXh/SetmOD8ZTuYTsIi0ovgu9KInXF7rFlUS
SOZagCi0YQxYaGCjYCb4S2Q40dfN7Dbs9hFap5MMaROlqzzPmibKRjxc2AlBttdU4dgph5zp8fop
Kwks/AETaR6/23uoBSROHbK6SqsaHUO56cYS6D9FYad2hEthM6X4cVAiOrislk8WaSRfcYsroYpk
t+4mXiMDA01yDZXETkxARKfYy2PzbHC0ehEC0d+PBe6nwiq8nh0Qm33XoBXSdEK1I6D+55q3TQS4
6MfCLIQm81ns0sWdlNVnZjj+U9mxYIzU8Ir3ovuBBm497ODJBq+LxIHjlnPgSzrtMDxzJFCb3//b
FXYvfs6ti7wieKgEKPthW8CCmxhzM0chCzv1R8YRxz8+l/FKZL6io1T6o7S5+bfyBXkSJgDGE3em
ic7e8ruu6tmWNS8wzLCuddnmoNTpegqr/xrQrReTc8U2d8OP042EHle6/2cT+stORj5z/0aIudq2
9buFbesZQCmm6jcH/1C8RruPs+gNe7jT2WwSdfvgkZcCDAvElWgLdK8Zi6f1kDHxNWlhezRvY2Qg
Vq2fLH7kS1gWh2areOPsREtdwI3LVc+MOJYfOVFLPYZXl4eEBsOTC9tZqg/XegHpWqlLD9A2KxbC
AapfgI5Nw83NxrvHPdp1pFfzq+u9gPYv8Xp2FBI4iP4Lmw7SCAXi/Mh2VaEKNe00F6aUACX9mv5p
DKvsLsbJ2NQBi+wP6BXd0TA6ZuxjV/NmJ9rbHBdNxrplxwKhPCmEgEUdF3KVo985BU6L1IAIU8Mj
cuvHxNmW+ge4NIz0ezqcou9Q0RKcRzhrbY1dEaEu8JXB44kNmr9Wfw8dXTZKQmu/y71cybG8umhp
sMdcc9sENnTeVAYBiT8rrY8hL53j+i78AQe7xDEc2M7PQH3Gib58vHhGJK4oIAaxp7KYKCDaPgyO
RYQm23jyAOw4mc53qySt2o7++/d6q6ke5R2CPx6p4+hZqPZvyC4w86qQqOFNjhriJEpVYa2OhERj
tr+OQ5GI8C2cfKI7jJoC543NOslouA1ZVHbjNJ8nqBqSZlp8xD+pZERyxylXFYjIktKlKkD0YXue
V+sRUjcsuIwq7imiQndNo1wjVYgIs2In8UCyK+ANgiFXKB3UutQn2OHz8PhlSiQfp/tWYfnhME3p
E5YBervX9vukQXtpS8GMts9jKUvLzaCF53WLc2+oSFAWY+7m3itfymAjL8KEcL9499W3IMH7Zl92
YQO97ZEH90bkQw7Pxh1zq8Zgn3QDZ5tqL3ciibRVVTeqkEdURDRPgH16ap33GULgyFVKQm8D5ser
TS19WZsUbNrA8sdV80U5240omuloOEQM3v/rW8aefUa+/LHU+DaSiolXXKTKA6hW+mEaGgAi6lzC
wvMzCASuqiNzD/0hGHGG5bodDT1v0/WIH12fSo21aSeTw7vIMgxUiQEs4ZVWv97+qtWxQfYI7DHe
pEN/iEyjG2eo73BzKZsz6eD7qgpaXHFMcg/7mp43nyRQBewvSjfDEN72sfhq+GpdUTua6Mbb2hgi
xuWj0vo5fR3yQC77na5QOfyfh6RrwFeyo/C6CadRROP/voaO6GuoKIijXEEv2gnwNVA3reXm9qKx
B/EZeSg4BV19xYCp9BS9DwVjWVbu1Ba5mC3jo7QVD7uIlVY2+1x7F7XrX13vjqJtH74t/RwtR1N1
Wvyj/31CghN0aj8RYOQuTidNNqUGKmiOrNgc8vfaLey4pU217Q6Th1IvRSTTOIvfqvcpdTo8XfZg
/+MPButLXBlCZM1YIkuvz+i4AlnIIrR0+euqs0aFWIdYSOFeYnumhsAEa43Z+6E4sDRaf4Ln/ZpH
JJwP3gj52ntf0A57eUo1JoiLB6dBqW4DFErRmd1AUCPrUcaMwjRy6thnyBjncz2zpg+AoxZkDFYs
+E+DGMVg9lkIsDsyPs4vrUtsrvn8rYR7lAEZNIKCuY3VMymEkxZObVznlezpKIsYlAFgvJPPgsoe
v7cIVMr+5YU7s7rlfiNf1h1vck02GDHcjqlM0MvuTJOHc4OCSGkPwSTR+p5A+G9x4DItKtDVMI1U
263X9PlzJdjaE32DpwYguN/PpgcScdiyPT5+FS9/thY0cGXIqzR3FfsvoGhGwDCxEtS1KcBP3jrv
QXZj5Vbs96IM8z/Gx8fA/oZzutrj7ctvUV9f3Qn46TrlTvHGP/UR8Fx1th3fHEAn5mxgDlGzn91u
k8pdtyXqV7JIwfGVrm4yV3IdPEGcs5DHc+Y9Wm4vvFZMd9F+9LEjddihs8WqkVGRS49Yz7fOx9wH
nizFSKNdwz/1uaJhi+ynrNSx0lncA2JOM7IwAJDVVUbMTb5ahajnSbjKk7Q0pm5M2uhUmbiIbIMj
gOjLqG7QeGEimMPVDIPfL5T/Y9kA01DAqJGu/eC/p7+fHf1N237SgaZbScBBZ637RMOfEZEudbUp
FxmfY5yFHA4DyIMDahR17kcW/CALWqYqWwtBMH0ANTqq9bTfsh2alKQvrs7KnPV2c1OQSSnHLxBE
7zfEUnrcJniyaNT8UMyz3/lqbYzZbQh6/UN/e1uknd1Tx2YgiQk8Li1mSsE5EK5aGlOVANR7Iz41
41mcYrevSJF0EtNW98/+kFte0pLKHMzUMHvP5Q18wsect4fRAhzIRTsl2Ow7bil0AN8bLHWAh1R8
D3UUxTILTJH1yQrABWbeloWURUFJIXjJA8cujkcITKFTuuU2F77DOqK2LgKYBPMOrDQaNrrjYw+L
yivBc/6AaHyHj8rQCNCk+BJHuVQK9AR3T2pPJD+saIpa7I8fWMp9OHiNUw8rdgaqylvigiuEVzMS
ahbpIOZaTLzjUtYCuwXt7Ly2c3TQml5PdE+n6WHbHef2MvbLaUNK6hPQ94deXaMIhY5Z4pnu4tU/
sp1+yu+xgrolH4NT5CcSITfju1Q6Ifz0WuR29upLjCrdV00q9up7If2Xcu1UUcaRKIvUoyyBU3xs
g7+ygyfMbVQCUXdTrazAVFZrKlJf7ZbJUVgmEJMIxvNUohRzN/kZulTCab7h7rbc5KG2Snz/Bws7
slaVeuZB1iXn4W7JB464uVJjHOgyW1mKhAlYg4QDUKnWnAIT3bT/2CctEBEccBkM1VqpknfTCgIv
1mc8bUU/kUoo98xFSnlIMzx9xXMoPxG1bmL3lEEI8L7JaQkhbEXhjVc2fGbyIXaZUUIMdu9tSOdG
12yNuvpurO2N3/TkFhf7C7JNHD77ibrbb+cZZPMUUMTnL8aA7vxwg5xhkScTp8StrxBhKmD1Zldz
9DZpqRFprbO6yy6ALdUaUHq+QunTNmZvuE1MS9XZ2EV7gMIV+NRg5LLeG9Wiv46s1VmShSYIpGHn
njKS9wDzib2cFHsSqCXYyJvFqT5rdzX1sND5FIiLthfWzhlC/pw/Alt6TvkWIg+Z7yT9j6ZiyM6+
G5PHQAuvAi8ckWg62JyEYqROHr4I2/rsGnsTFWZO3yxtMMRTwrKGXlPB1VUDMXGwkG+T7xaPkPy3
EvbTu3GfF+l1BqxxcRI2cx8la2uGRH6S5MMA/EcR9w5kO7Szeo1oZ90i+WWkBUhykBV0i2kyYFhB
LnS3Hly97bgFgkb944O2BrTBcvD6OsVOdMQd8XLn6SbVbcnJqQwUUawxXtZT8LIYVjouFdsztCsr
tKCzp5PCKh+wvk+645Nse5LinubboYzybrjL7aaLLdZ+tBWumxw1DKgyfMizcPgcpzuDqRtIlJLP
mlkWUMuLNpR28Rfk8qxGbXkhdDB8xyfWEa5MxYSOWda08VvfK6QP63hTBjnVOZkf/gDLh+KdQ9Vs
HA/hKuDaUEYO7e4lB3qZ0E14BVyoxkAgtDmgChcQLZ6BqAmtU6rsLNSNVUbJUTiqzRQTC1t5lqQl
D8A56+6LRrPcvaCFaPb+lDtNyO8e5BVXOtdIGIwKqPCBI6yG9GDc2Mn94vDKdVc8/FW0cMIohbGD
h8HK61yQ1x0pwjBYjEKfpXIhQ7CJsCtCNnewOby1MvIuov1xQfyuZ0R1rlUKjAYUwLtM+HiKBPVA
1XYwDpNMPsbKX8kJ0km5rjf8duGdHE+bTw2bKqvJLTKeWQ7aXpJGB19RasBd8vYvJmn0P0Emix2f
L0c2bU5MHb4FhttEd+IrNRqyODs24nGAfOdBHa96iTfuEyYZn586kEGiVrTnBOcfLO5eB9fH10S0
X2gmrKHYWpNrjCtArHu73qZYM6N2Jp7YA6T3ifcp48oi3B6ou7p5ekps3JYK3Ia90eblsNsIZGXq
Qv/DfrPOCKEBD0R2R0iZ4r7QyoVml6WEs1lhHR5zkJGn5W6Xk0ioriSnbJbCT8d3syMmoCgxgHLJ
L08+dneg2o7AzYxUcaZL8D3y26QULiYzoXQ8vLlB1sq/1KkLggRP7OV+5ydrIhY1MV6NNEnyfYAD
4wnFL6fNfzZ1tEGhBxsOysVGqWmStIiQ2h+FNYAA72+t3+EWJMpJLKmwUmlehJIXVVq9PSb8rIjU
ZH44g3Ujal7nmzfYK2+4HUBQ18lz0MANiGD8m9BGO9dL/YsT9xryeWGl0G6IWQ6UhA6PR15Abv/5
e4IXePeJLaJGezhynZhEbhsjKEUfnr6H7dWfM2zyRM0Ve9hFiRv+9SrePvBD/tLmF0YOzmvnnPxT
ffhFP+moecF/gN7Y1nR3Nic+MX7WwdyW/PNTwi4fTYs8mUZtjSTcAKvl+rmGlM3FHDCOPLH1IN/H
4YYg3XeKtuR4jbaIgijvpgDG7/hXnz0IH78nmhiJS1rpQoSn7zOU4UmCh7PY1VpIXB2mHsPDzUo+
LlMaNGpcY4kt6qT5y6+t05RRduH5JDmlmlVVvDiLsSnFseK3k7/JkmkbVYIaL6gFLH4M9wREv28r
D/FYVeSMTHHtu5GY42nJBOnvCCiF9Rm/H94MpWwoKXiEhAhi5XIGEEx22trROON+ygbC7kN0DvGp
2e3NvjtHM1jqE6LFOs5oxLR3OSPGH6cXgzUVdd5t9D/qRClc5+WBJGZVSAd5wLo2JkQ6ujJD1GHt
xMz5xXZ/zkX/4SWsY0sCGKaE4TJvl/tMQfQ0L3tEHvTSpMK3TI+gR4dBL7MAY/boQq0LSIT1pQRk
SH5pzqJtLk6KxFlwAMDkUhhJl27jKD3ROq6pzsOPriU9vdgoF9PljxDNSYYqcePVH5T9rXzesuvM
brR/4kU6npPaMwZNrdpRUo0Yns11s44eJMXs1eLJx0KZyv3O3wlITphXTvarnZ35sRr4h03Frpu1
tSTS4+/UTlnijo7/2lr/Eq9ln3BLSkQObWuyp6mu1nHytK2zj/uY0Rd5Nz4QineLrj+DQWx3b0zL
xZhS8ZblYX7VUL/jWeYRB6zuAib2S1h4Rgd3BM0C2IaRDz4aGvwXLII0LMApMuFNT+tBoCN9W7N8
qclNjHAxuUKnWjm6n1hcFshp92V4HNzWrEvvVb0u/HSQE+VHRhiDMReKo+WgcL45cnT469VPRthr
6O7SfAXnCxECcx7x3YayZ4cb0RDYcQ6Te5lgIpe6ClrHTdfi3/yhVGRlpUNIYWVxps21lpA7JXjc
GnpoGwaOtSIRGmdwxm3dDrt1j3ArsnkmMy54z3bNgQ4B+vLRyRB3z1GutCpHrT4iOE0W4eJF7su8
yuqIW6qfUVmoPv3SyEl/BDfWoT4iByoqNwFyeZ8MY4L/ew9RAZckL9ZNxT1lF9bGo0NS3NzaaA9C
fnShhCZAl3Vdh9aF3ogBgHBH6qInzU+AsxtB9OBb0kD0BsAsvM+Aw8YS3n1mh+O4rqjO/twzceSQ
TdqBUlSlH76rL+lFTYJt/k2mB24ALM+cq+5nE7D5YsovnFdjXICw0SVvkL03OeqHOOAzXcshxvNB
fK8FcqzFeFNE3SauPPFiraLfe/N/4+6NM2xOSvhJVi5V5BQCLrxlzgW6p8pOoHAXrebDyW4D2Bn2
BEekHuz8AdvTJgZDp0cBWhMpIGagl6dI5Zeo9TjdoMKDC3LxLjuoYrON9LIJ5Q1Rno+NQbMyqK/z
E+WXdwZOfPm+hD7puDzGEWikd2E+JoxKxIv33DhBsYrOWgoBBMl19TqHHA8RO4YTjiw0lDasDXFr
TQUAsaJ3mGG3n/CzPhJh25v6m3ry/eDk+litiA8mw/6YYgDMNjBgdxkpoDWvINn71pJy2gJIHf7B
WicBlSYvP/mNKrieeQXFXjNqyU12/0xTW+i0U7ztvKzISigoz3msJRqv4jgdJS3u67LbEzdFZm41
u2+bb/KGAifejrPnNJSYtmPXLQPIaWyulRbLwsCOVkSfqXTUriO4eNwfTfgotdBX5Wze4idf3mL5
P4z4TYTEr+x/nu2TKRC4SuVFDJWp4Yz7XVXqzzMZ/zO+Latdi0+VmnW8A6x+FDa8VLs0OMHULknc
PzmUtNiax7ASOnZDX2eTLzvNEEQD9ZCaXyA1jqc2XFjZYjjUaA1mk3wvW1qtB20GAZuWJCaBKo4c
iUOqaaRV4SpDM0jxVJPYheQo4OGvZQKkXUO0jspTK/ZxdZ16WxHvQB8zZ1r7PBfn0FrFX/4vkwI2
77rtuL60zJW9EVISlIZzoYJmMgBZvZAgfqaiJMqUcTjRGq2EOImB6QZzpyX+QfirtyLpBNnUIdUY
Ppwm8uK1yNEyTlm8kYn+/ZUDZSa6YoogUFS1H0hGmGWhNz+G/cGF0bqSUVQdko9FSXcKYAcw/8HS
YC4NwrvaZ8RSDgc9f/zjDUtE/9v9KO9xC1ck/dxM812CAqqagiemEuiH29O7M/s8jhiIlk9gvGBG
mcPoyBImmNB12e+aEaEdGPwRNFIYoVMNve8lqMMd8x8iAgMW3A38hQfroZmqD7/sMWzHJAVI+V1N
K7Bh9CxeQUtDk786Y3u+jBgVgFGClvHXn+irbkt91DI7R67jwgn8Rj7tJXDiNJtCqmFmN5+pWHRE
2v25geg5mZSz2XIo+fMRjrb6KEw7DTXEY+7qeHBEz7zQjvQoN+jY21fBbLGA4fPC0bLpmBXM/R1m
Kr7bZVxhUqBCMCi00rZpAMkKFSHGi9PaInSQVVZH5XnkxbUiSmZE3ijpY9nrYyjSucslmdNuPtrq
kAic3aB552YXivRsgAHa29uQKAeTlKem2e2joB4SQHTbwx/T8+etNKUal2QE2TKDVuDCjUKZ5d5f
Hno3M81XAZvmAIAlEPxxy3Ke/mgPmJlGGd9EHKRE/FHNBEdYBjxDTcSjSz2mNdJF799D8k2MutNK
1bYFdzKkoZ0TYenTLnUsuZo473jSuXVsdCsLWvnN36jZUT6p6t9LtqeOpMMgpEA7vMBrVtQUuP9U
qEe8KbgAxeoVwKxtOCzEievEF6zT6fMUjSOLWj2BWm02/TXBw8XeczvuWy5eJq57aWouGtZ0nTzh
6207qNSFAlwWf5cHaj4pi/BeHAlUwb3ylhCnElJjfiIylqg+VfJfFTIJHhjmBtr3me6j/LnhrHXl
OBspJ85sWW4+Mxw2Xt+asVoMzfX58/5hPf64UHEbuAAulo99sx39Fl6F3xFPtXRifoInxBeo0kKV
Rw6DCBPqFIlYgiWBo8umz+RA78CG6GT3ujZe5UJnG8ep9fPZNIwAbiQx+fxA3Oes/k4qLmGcQAsl
VOPpJXlygKjuoZHa73DPxGMHkPw0Y4BO1ePZXyo6ijkSEuWJUZV8hgS5U7xz6vYcwt1uhcPaD22g
eIqjzNZ5yyAYKY+F+5jxQAqbzXV8N7iJ6h8vXjEk4Odcen11nzTzUHq5ESnOcpKD+NnqyOtOTQpb
KjebCtxepfiZ3ynh2620k6RfhfMg8eTRe8NuJ4JVbgwM9pV5V4JHYkkoq+1Cz5HdwYiYhDKEYx12
NYtSf0Xewmza2mDSbnHOdmJ3DNiIlJEBpT+azqgibdj2PbSFUIyY9crJZ2GeiL/pkj5xq5SaXZO5
bYTyPqlpPjxqeaEDN6kCShjdunasZ+BBtqsxKM+MfHZRcqkv+cdkIepmUmF9nd3myyGMs18s/klE
Hp/m+0Rk9/AgSwF6XSOAu9PLpOcGQIPix+wGrQM4Oz06h3WYO8gxKzmwp98QwV+RhzsuxZneRSAk
5qTJmiH/L2lj0FRHcHkVSp7wISye9TSxV04pjZ4xuZck/YJogs2fJQZV0K+67GRNgMDVGaGrSRuK
tgkpsGl78rJ3U0Pf4l/bp7I48ssMkwPu9suwyM5Om90M10JCUb3Q7iQGeqFqs+lFPJsHxXJ7JX7S
A1DxUnhyvuSpiybyfFfN3legslA8WCJeSx5XXHUWBzuhudJ1v6Hg8Af5PqMiSwOTX/0GXy44oROa
kZZLowo4oQBWQVgUPYYotzhUAncgRc19erbg89Ht6BO5+GamNKC6jyV8ijymkA8KZlzN/TJbaE6m
q+OC3nraX/IOAq1SF1lh78M5nsDJ82tnRXy7w2vbURWh4fuiJTCwwUJ0p8t63d+dqWag7xLwznXa
uw947uMBpaylCC4KKIaRtabqq2U4H2Ow3HziUxoRcjATrj6gEQBABzWYnIgJ10lmBiy3q8XDswTv
ffwF9ABp0DcMWeuflJ4ZdgvNII08rguD7a0YYL31ZIKEMItEoIVah04HdVg5kXqpDe8cZX9ehVq2
7xU9umbk2a8zzRgHtl8U+f98A4BBEFTsOPJCh27Cr/5iusrIy0hGE38OhyYvRarQP+rElLyKlpi/
34oQkrJst3zU3+tV+HQULzSz/+EGpOS8yU+OKR3rO9XhTeCpG/P48b8Y28liaG/QRfEbaAk0IEeM
FYyhXmEWmhVr6t5e/GzymML8ETWuD/S0IcEW7L+aMCMRC22oqF4yi5YCW1Bf+zN46o+eKK3r9c3C
8sJWw2T4LdwwiKqixiCrb+iYI2MKYIgJHv2wtOy5xIdet1U0mLa4OhRNY1FyTuGaAepUrlIQmnQF
vZQILzgoiUxTA2cY1roZvYMz4sg44q4AXt0dVjqZRzc+lLE8rX6QIzrYOofrrkUVyxJbnJWHjzAS
bWfIPt5ISdOzH1RgXgAvhOvbNSmNcy+/MLlrxtNkDv5kgspFjpMF0TE02whNOwUiENsWs19GGtip
xUs7BDhQu6DWGG31plZZi+iwm8iklAQyIwnMXpSA9uKRov5lAg+2zPxoEnV+5MoSBBV0NcwxkFQa
QBYjbJCVk03aj5w0yRMbAGdEzEfdrB7Ee1rcSNcw2Y6resxW2ARd9ajKB6tTmNVndiE/0XJSR0qN
wFVt4Te6pKTKFMVUGkJmYFTImBXnz13LmpGxUu+gUIwIIjVyCCb8DZO64KEjS/o89oBPZgYnlKOF
X0TBT9LlrWqPejF1EmDHHVriX7mpovWtwem0C4fw85mNc0TkdqA5CkpXC/FfK8cPg4z/PBOEnF9W
CmSodkSO/yhgxeLS+mL7eT6lUfI+lfUurHoQMHau65hikTvg7ci7RU5j7eyttred8wzEjRZRtaeC
bN84CRvGij5XCHIZehHHFB0TxMMvhJqt5u20TELhrKSWJQPYFI7VNs76hfV3FqUTjDtUO7qm+cwi
x8TVNbUgI3dk+CleaiEhcJKKQY2OoZ0DVuhTtAXIs842TXxkgujsgJ52cRO/7Nhe3EUGSSBd/C2g
3a3OFfnDSNHC2dFMcFmboYbA6D8eI7f+I25rOFvYQ/sJew5Olp+L4FjKHlzR6f7zR/dKxl3us7hF
HjEcvMexY+AOtVe/gknuqueCxzVdBDw7oBgO9czV9DNquXKOawr7DsEQTXrkrDao/0BWi1//tCrF
z1pJEAR+XVw2OOS/2mijogy5Rd/nwBKH69bQW19GcutfduqV0RO2b59bOVrwfQdop/qAyJXMubV5
dORYII3ePL1T9T04iW0XaYxgLYjQTK7PwfQKeCP5a5+8XAzR+XQrGD1m4c3NBMGwBYb9A5yyZQpZ
AY6doHN8JXsBUHC7VGCmfJdv8eEM4ie/nuMMEvuUDUyaTKx0MnbyvfByQBUFS4Rqky/2EA63+Kav
E1FQUJH0X+Ti2+IT8DaL42lHK2w0Bn4MOPwOPo6VpeVRw2+PMYpfHIxFsLeGoAOtkSzz49iX2546
vC0KPBdxTLEIBXgPjRb/sUQr1S9NM8NTli6JinY4Wz1k0vdRFphwOOTBJ0nmFJCq+KiyLcFzECgn
RJRd8wgmR+3keP3GOh0DIu/UaDcHYZHUUdksb6TKTcgervwPcrQHQRitCkhkoS9niepAb0Lvv4zy
9KVDDEMnnGu/XMOA0HsoKkw1cLTvSUetnXgjhZy/kE+dVBVteV3b0YRzNMWuyovVCENpSkao5NkU
vI4IBs/Z/AlCe/Tq344tv41J/3PP3XDMAydIh0Hz6SndfCucC0tr7UI7BsGcA5h1sTgGkHvDFvKp
ZHJQLN/BGSlEJbF6eeKWm7sPEYNZUKaagHVE2fB1r/Z8ba0mDGrDln6mw4CKQM2Tne3CZ6vnziZn
KNSZ4JTV8LOPE9OjCjnBXBUYsuyR0IqoBL6uYYgJ4eOt0bDHVCbCIdEqYmIJTt6ofJVXD0afcYYq
y1NLz5v5fdz3PlBnyIiJtneU1vfnkoW6pst/t9P+ftn9jp4pqIIkA+HnLbYG+mlpPbbvHug8sGvp
KZqTeROjyF8JAQc2vUFqU/23BsZ+heoyFMDdOGC8EtfVG0NwZQZ+DGd/ndtqcCzz0F3tAEnZVFc2
YzpIj1MrJvo6F+ThhqkMiQxazje/f6Pf2Aq2nVa7siwiyFb/clYFawnb+cSIlNJi2Am6mfwd4trp
GyQsPCm6Ib4o6Y9vz5FeiLWjykmMCc0Wqc2NJA67sXf7roFPBnTXRGNWRpBUnnb4YZBbMTqT2JCk
2Rg/nbgy/bfxJWVt2lsi8OwjXKxQWSFz3Qlnz1PTk7zVXzAiUAjetG17xxPbkXikQLkayJZ9iSVn
IAv+g7aRh9MlsSU8kQoCOX7aC3f3UeT7uy1Ao+GeD9lqj+bhx/llDX3XBHW1Yk2z4YtFKeL0qimB
OgEdEW2kJMO9n+oixyMhsNeRbhDDUijjGl1W2XUA8oVvUGqrTkEEZ5ENt9rU3/EjjyJgs+rJFQxL
nOw0vlnpvCwCl5ViDTq2Y/Q0fe1awSWyfBuVnwM6+g/EA8gQwlYbIy9rBpPbfpxQFdNB9pyc/P5V
nYbHWCRoxJfOZ632hekS6vBs1ryOQqSt90Tei3wwwmMQgQHnNZcoV88ASFgr7zYntMoWwcvyod16
ZoAIzYVK9z3vAIxyKAujY0pTxqx6b2ijojHqOd73qvw961nph5nvKfyAyWotBg0t7k7n8+ohnfmI
npwETDjyzfVqbWRKBrNjZYJl1sv3kgwnB/yW0DnTNSrAVK0+0Z1iKqOaA/fI0ZLSE5S2GiuC4hAx
sr6CsGDJboAo45Cqo35Gauy4HHLqrbu5mb7i+GeL6JgIoEbVTMYc34ueXmk2YmdjXh9VuAW3pB/V
hYJFvtraqWeXsNYxdWZeDIIhcE0vvIjDFfedBufX4KEGMuuoZG49U0bZ/UOZTtWe83pHJuQhVRG3
QzHGnZMQF3FOTtrIXTeNNE2S8xtav+dWF5ANfAjzV0ncMBhFTBji9phCpbJzqWUoh8PgtuxtPsAl
iOdUaBQYqZ0JS5kIn6vUFdbFZrg08o2pahfgZFuiXFcn03rhLHNtZgNclw7kWntWFdZqlsZsTMf5
wY+hoJtyDxqR/y5uPH98W0+bo8xXeQ34UP18eYsMfShYG8tnAOl5jQ2cBN20o/qUpQtv43cRlWDb
HCMI2uZQSDtZZh26jSo3IvugnbYNi88+yOVFKPbNNnKWtAnfCkq/dkeO/f45EBGQxmAe0ywHesAZ
1GRZljZERJiv23XRgh7Bh1CPHlHB7BdQUGn77ipYjFnJc76LYIbeFzLLQQnpW/9jjRniOQ53MOzO
DRamobMFxbEMR2iLB1L0idB4HCYSzXWicVPATQpAmJb2pQQsB5Igio+wVNVcgsXNauGyir5QcRjI
+tgpXafBFeDAhLEXn4/GSViqRzg6NOb75BFRv8gV/Kk699o/OZnzDgyhUBhN8grchpTLi2PYdICw
MxA+Eaz85Mcrz+SqOor6wceDUjWjNZ0bGascPc57NbAa5nrpPVQt87xoo+cR/UN+Kn26x0lfdsoL
Tnb20eOCHNRGPyrQeFn/UEorl8xTpBAPzaEaH2yFwx6/4uXJmQezmHRvqSf6JAK9bM/YkjdDhfcC
B9YGsnmui5BFcxS54ypv0EuEYHd6ZTC9cE4xoz6S8tB1SAJ8BuNAlS+NeoQ/BS4DIP27yOgK4lvW
j2EIOa9aOWkB0D4ngc8LJsutcDpXwGG7/cFTO3Ko5u2qyJylN1mqEEav4lxlXXKb3IK11PUfC8Gs
JXaoHRHpk6LZXrPjnCBmtm/9I0WfGsjas+doOi3Z2YftfCZDhUE+uEDMqdbOKNCMJZ8w/CHKCH7m
nHU6dAOA+YoJPHqn1j+W8K5MC9rd6wYuQyPMutrKX1UrZoETtSeMRArlBR0gGHUeh7VmU+nbIIFi
8G1SXgaIX7BG3PEa8jN8v4ux+hxkDMmToHk5a3GTN1DLyeMCMr8OVLKKImerMdRHmK6N3bgO0hYr
TvDuCeqSv4YumgFUwOCYZ1SAYReEHhDqx49ovUZZlq1zl9zPuxoODc17DS758nZNMAhqOtkaE+ce
maaIF67NSO1RKyzADFOr389FrlZFK7W1fYRpRH5+dAbbwrQCy/87gWLFeKww7BAybPzScBWrK4f8
yGdgPgmhCN2Uom5ELy6S/fHHUH35hGczxQIkQeOaPhpo6UuwuvBBjkE23WtPsHvy3x5sovwi+lgy
tcTDidFdddQ0cjgT+JFtB9TNTGW7cQy51FoU4wGxS4ri90X9E6cKbG/7K7B+hqgRtdf8oTZ/wGSl
5TIiARz+dXj/gL1jVycBkaioGgzL5wnvkpDDDief2zTeCapVjaA4rtRdF3KahJ72K4+0P6wV7UPo
XlRC1FpVDjqF6p5zgfZXitpKkGKKfv2/8DYbMaFv2GFRkRSsVPRnuDjA2+AEgnW6ExxP5vDWm3Tz
bXpcKgeSBqsHQmG3uwzPrA5yByDzrdojawKESVfW4QhOfsB28dLIQTt1xi/DRWihnDu769uY1QBY
hG/LUm9xW0ESKqNjZjx7wK4tbpe5zGqnWyPtE5rvPE2OTDGtIbjPAXzP8qOEj1P1tiDHhyYejjbf
ztVl19oDUN1nD+ZrpffPD3kA6TYOtXd53T3VAq2FmbTpAGE5IyEy+n5quaAYqJaiT8SGsqL/nzvu
MA3EfWKFKowpd00By4YP5YetoWQuI3l3wetONHmixz1ykgCuLbJPKADQfSbmBCGIlOFUjYbI/bvk
PPp9oY6Ix/9Crqj5DGa2ByIw2Q9FHCzx2tDCoSDB7+MhH7PGqM0H5Lww+xWZxrmDO65DPORD8wRa
mhrKLSiZCKHRj48RZmaOLN50SksDDC7Gm+XbjISuS2eR5TAnhYt4FD3ihvbeAMql5bMSIK977HRj
1oS8Rrn4i1J9Z2wgcj/SSYYOvpHXbJ3k1B+e8c34Nfl2ujArX9YGoKB9cVkVmnmdTVWZdlKN64rf
i6rpJU2N2IDd1yjbvdGuyppQFJ5P92O3zL9ODxw+14WNK3OlvRzBBi0in1nImb2CBY/LN3yJ9PFb
ch2sXoIeiOIUM5oW4onPu1FLb1SaWvQak8vWQo4/hM3vwgw+rkjO1KGmVAy1kMKiwzDq73zcHIIc
hX4CGunCmvrWIoHrTxT96HAngYKaT5YsxndK0kn/FgMy/Q1Gh9NDdY8365IIPyUl9NZXwtleH1k2
Fx/u7hUtOc/Me6IEXDAsy4TnTrWU1TSG1lkBOxvgT0iHD03RJ6vEXDpDyKzNbXzXdttygeP78qUj
6spa6yPNmqh2Op3M6ZVWxr8gRgu6mwJERGaUVLCAmAVebUiHXfw76Q5lHaJiH/ecUA0+apnHwk8b
it7EQXl8j9WbWmRpcEK411kmXxI7IXgjD3H53GKB02ukO/7d2/jRPz81zpXxcqCpBL8S/waSEIXi
7rO8heOcPtcL3GeFq1h9nJ7Ttpa16/zOO+0RVFbFHuth8w4IDsuPotu5WzTALkWkAZzE6nYau0Gp
NnU+ykY/seO32pdyRwPxeZDjtyI3hpUR4FYBuU2kbGaUCHeBdDwpLGcsHrjkGdB+FGkbt7nUQavX
e87Gg6kyBm79A/O+zd2xfrJ8t5ZvckIvLpV/lroGrrjczr0xoum4h7M6C/rm2uPKNr7phteugiGl
LVpVbEPOZJEWes4Hl3GcygWzigEgObP6C76BIr9PXkC0h9nLDgqPZoYWK9TLjrr4y0s3htUEGVRj
UMD9F4m5q5TH+FNt14GJb6Aq0HXjUImZuKWgCMc/Y0NCA7cTzbiq8OONFqYHvoepZ9ipYHZgzMf+
PZS5t1aWZJ/jyOgagzLciUZSH3hd5nhiyZApdgKieyQmWw2iPhf0PEYtvw9Sm2wdYs8rv29a4ANy
8pRE2vrK1g4v2vqGQRvhda/2s2O1YW3nP4Qb4bPkiJ4TxkulBZpqujzLKgW0O3KG2o0YNTrdIX5I
zuB48zMV5yTCzCENFmIvywyiAgVynzBpfryLB+Ya0h0Ojy1/4QFOxT6D5JtMRmrGL6pWtcJ4rJ1l
jsMEWEOt1ugyidAZy9ElRuGzLwa85MIPV3SExOkXWgV08kSsi1h83eUAaYjIlZ1qi1xwFgDDmre5
JcbRmiJyuT/hE0mGtENDqYfAVoXvwhpoDiQjBQGSFhwc1NLmUCbeUihriH480mDd1qO8swTJeHjE
EuZ3UUf6mvsEn3yz6ioTxNsitpPUs3h1DqkbdyxEc8hRnHjK1vGW6oB8zAxG02sCQo0eB1TAI+Oy
pquXyrRN4hU6HvpTrnjch4J/7xTErbPATpqwxIfIwpA1Qjq3g6h5zCimRdDhL/+ku9K69QAGaGgG
i76Szkoi21D/WggTHrFlfSnys/7pBrK+Ch661zBPneP1YqZazH4LQhtc3gpVFdoROFLdFllfzLa/
lNGgtlZc8oEnuxny1pJmnHhfdHomEzebYcQaYLl47VW4sRWl1PWP4qHNjsUodqNxXNwa1xDfDRkS
xH9sVJKVM/Hc95eXP3EJIp8wUjjEuI4FJTG2o8QwTPEaqSVH4ywCQDqPbrzOWQnscdjJK7QQ/aTP
Yo4glvgu48J/JdarHFV9IhUCgQpwUB7QKYRKQC295nSraHV8t/KbnxcgvmmD+VpZ+st8c/08HLzy
6PZKOxqAr5rcGvBvyXh2sMHxQyJiOxJZXYASrmOr2/foEliY1uLFLcmkVDxp6i1UmRsav7gZyvti
og/N42W8SXo12MxGYxzDXFeU7J2wY4fCYacYijH79G+YF/kUMhKytNxHSFzVgwgyHKnYQtjZnc32
IWtLvcFzSGrRr6G6OpnEtvqDXSBgdCPGszkPeXVSHdwJDEtPROcAQRD0MsL+kTu4bo8iiZazn2kl
KtoorBXFlWS2TdalHorplqJc7MM0ofIWRHlcj/x1g3ch9DW7Td2lMZP/66JM7EphLt1m5Y11EtbX
XZu1aH11zMrXrr8Kcv7XiDE6UH8sWx4DMrdhCCRrgjIh/88cz+u9o8psPCC5xMiSxmqp7QQD5VSI
4QINWTz9Rm00Jg7NN4r3Mm5/LPYljnC7UeFmbMHa1oQtoMsjxBond5abv4o2AYQvxGluEkmZ2L+d
ByL35qsyQ8Svb5j9wXqjFLp1t0bHKPDCBBRNR7ops22p4FW2kRvNBWCTtlXgvM+UKKwr9DJcqLy8
IcQTsTLkqSs4wvkPxMf94blzzsqjEEKI4Ifi0aSjh0tmUF20TTvbcBdLC3aw6Ixpld472hkwwjHE
7hpkiFr2nHIwEEvnkKg8ECZA5iS/XzkslbiksNIdBR93BxvzPEaxU9SkDX7X/hX2jMcKBO5GVOlY
pMV7fS8yRErlWtwfmlUi3GlN+/cbuum0fc/6Hi5r15nIpmRcVWFRWtkiEO4Yjo/08ry1ia2KcTaM
9MX0Vp28cuAeTEkKT0EQvQ7R5otmQ6O/7k/4MbHzvOoyNcbPXQrnbFHoUmBQ7TkEZT95eRGB/hJE
SBf2TR1YXNDfrEx4BYDmLWCt7Dyd+HHhFOAl7S7ZaVkXlvKspNsZJW1BPq1ciy3/5eFKdPcrnyu1
miPIyWbyEoECh7YnoDg+e+exV8aUpvsoowm3ZhtpOwpV93Er5gbxOSgr9+8PSw3Kv5awFqKPrT95
QVev0no9BBP5Z2FDJYRYv8/VI9aN2LQAzq0I5162W3e8oUYmh8h46yFPIAS4OcoTFg7jXxMPVWrj
zyyTrPz0IEpZ5wr8zl9rZVg8ZkZqsgvfEiFIq5b5spzRYMV26dD1m1X/SZp84JeZ4luyXeDXbnk8
XD6b53mDRthCKT4zjLnn7U5PN7G7R40Zb1t43WUIYINKbHDvK3ZgsxFdd4MLOx9FgRfRM8eI9yun
wBErwapo1T9MbS19kLfPQX1Iq6q4SxdNeLS/flT4b2SLWIc9H/ey8fRscR+/cpFUUr+1xjcgG/7n
q2I7OpLDCUuOJrAb+Dp5/koG//gQHH8lKx3DRSfFD6c4ZkYb7bl2UFnMX5PRLvy17ilMzbpGWPEl
e6ATLuhxplcFIQgo4duatJP+r1CXrq3thVUGi2PXKH/so6utmrj9G1SW7Ivi1JgUgaEf577GHshM
UL/ZH66MT+dnPrpiBt3Ch5lJ8sBcLnIGCS2HnnGC3O5/siaQLUA+BHgjAjF7K9ZxyyW7O9lFcb7M
a4GUwQPocvubFPFokmV0CgMflxa68s9M5ovP434aAK9BlL9JBSC5wlxVkVTLddNg05UFqm8xJyP5
+L/DGPK2TVRnMksJ59D6kD4ea9lz51GZtohCH50RzZ6m9btE+O9TbHxS5Uw2R0+WJOnu6aPb9yID
SgF7PL3AQIoWaZuh8OpCLvz6A67CV4tlUweFvFBlctVAqSZqj8p4NcX/0+RhODtxrYzdT/tyB7rn
/g21Ts1MQPcnpgMrqDOVlCF2y+I7EUZ3GcSmCTXdDhUROSHAiuCN2bNBGR8NDMA3YMMJOAnTTT4T
vNxdNSAlqzpgjjntPPBX7i+0XaxmveJEgnY9W8BM0Lp7fcuFgqmdeXhytaDBF0vhJmRTIfhIxcWw
idH84q08WQcO0gloL9be5dNLRhaVEjnHOlrvikF2mZDiqmRfR+oJfVJswuVnZ8gp2BRKcRSx7Wm3
5kjCTSJqt1Rx44zn7TEG/PGB50pSdXfJbObiQT5ZuqQnbEW+FT93o2+94RPEbyz4Gv+zwYhFGzqp
J/GRBm2HkErxqT35MnIbfVnpjloIdtDKUAQ+MpQJYZE20PAE6N9iXuO1JAMZM5SFWBp43IwDJgYc
Bv+6WPAq95TfztnxlyaFje2SInKfsJW4Z/qRvhUisVCZPKVRaC22ZOpumqEVK1OsgnKYTva411Ro
VDWPEW/6gYEz06rd3WNI4F72h2FdCWce1Z38sdbAScJn8/OK8NuZb8cCaXfD0oL1B4cdCuMkuHgz
tczac9aQDhdKJfXi15s+m9sHedAMmcWMQji2Th6HyVkGyLmbGMawXKaKuKcXILwjE0pL2VDvsfH6
GYAC45DWfixWpq3Ll3ayhw9tkvR7NkgN8Qouke3xJFs9jJ0cwXDwlUbofkZkHvjgIwtqEuAjq3xy
WxwkcZvaZ9fjPaHLjgNKn4iQBsjYDMSZC4zP6hy5PtKlYwOEGI/H7jF/9eUE0huX03Pkok4ehu88
6f3d38FV3ePqbhzcODJfTBBlZLx1aJfWkIdn6ajknnS3xy4eu2T8HuE/TgxtT69fRuI8kc9jkWZg
b/4Gk/P3CvY7GTkqd1cepCRV7ft54GEp31G0iGhIhexCMomDaBOtSekSHjyEcmu0cPs99GewKdAd
W1qCjRMwI4S+VU5R8ZXZIzeGApFl8nISZqI2yi76d2FVdh0JOxQULfpBlD/Fmpv3VkOKauhwjt5J
HTD/MJ0lWR4tS8gaoW0zH0fA+ppiySkj+ey9AaY1WjvQd/FXRV+gpa2SFQNgrRwLLcvHVciiRoCb
MPwUNI6zCqVTYKp27rHjHvnvjV4bgC99oNsFlCQj8cFSEyPE7FfwOtko5LDsDUE30/zID1e++d+K
8DVdeQvx7QQOhFdlAqtJ7S88cfz0nauseb4t7ViTc6ZTgIcfGPh302136r7N7WMtN71lO6a753OQ
GeY9AQDH6i5Prd9cKQCoYpn2hx8bhzxO5kYN+p7SKBSL4iyIj9TZBFvaNdBuiZX0RhhRb+MbWSuo
QTJECV+iF/7H13wY0rzSHvKLD2uYipNNFZCrW2cBAOi0uSpJhh81rI0NxjICvUjhvlQtWEmPtlrX
2nRECc/txteVvPQqcjQG0G7kaTX/+COr1KgEsJDH//AGH95AFDcwaf47FHE8h6erdz8mxtcxAhz/
YGlZIiwrEUL7Pb5oPM4wLSXN3rxcks+Y7Dv+IzJSXUu5vWkbh4BrcBS+AWhy6OCwztVp6xF9J2Mz
0qQvbARBuEodp/14eN652r2ZrWrEFWsslvISzq53N96v0QwILc57wEhr5odQE7QbCtVhVK36Mg/z
x2AkiW13byfxGnUdr1TVgBx6B3oPcjsqxJ+n9AFEj0MTMfDsP9Opr4gYDlsyvMcN+ELdjitj2l+v
y3p02jdsJ5hnRSzguNuAkQ9h9lv+i0ydtYdpDYzaAWg0YnGntuhuvPj/P07wssGt+B0xef4z8NCw
MYGKUGwxTHiFl6anbPHovDZu/Ou498jTU9iMdtVWAiYvhc1JLKnm5IFDVl8e48a8fhkR+bYJfzUJ
ka45Ti41kF70+k6kY3NZC3Nk4JVFIzG8kbx/3vE0rmTWrV1R0fGipXi+j+B0XzNMBlZTsAWkhLqN
SrRyQkDSQpb04VWbvTJzAM2nJQsxK2qOcHOETigdp3bkE+WpCunw1nwFeuG8cVLh+dvIwkWr5JVP
okhnaV5nhhp0O0BtXw1guYmjbDbhqPoJiizShjCGEXhXxR2jYqL5diGUJj9D9YWpyWtCVJ7RPI+u
QCP7gRxIdLRqklZj2C7mN29Nux/q2QWmvyKH+EOQ6X+8m/61LDtFeZ7epoyocbqcO5VDZ0YNq4EO
EY4Y3L8ZFkzL8heF2s1XNTnTd4OFB4VcXyLslxcokU435h67ErmKlRsl07ZQLmyMu9R5BuboqiUd
M0CRef1GaeUJkEIZTw5/ijr/HCTVL1DSIGwCrrAQvo0v63gyKxWpWsNQH19EamUKLZAZlgyP9bWO
RZazGKBGxjpNUcdPfYf5Q9Pu91Vlr7ijZQ4kGV62aBWLTWzrDfY3mDBPZn5otUndZUUsWR6sWhbp
GJpmpUYXOACD9cUvWO2vyQ51AVc2DJ1HG4GBDcgHPtkkYu2FU0/ozwMAjn3+otAYXxHWHhpzu2iF
n5GtWiIdlsHRJvWkqLzxSwunb5CNL2WNzvrOEvQCKlCuNFbz755MDrIhdBPBytVTZkX3gCxS1uHa
yNylSnaNE3e7PiQB+0qqXG91wE9Gp5FhK3q8C1i+xmcpX5dBR4rFiilQ1elUSTBejlObuIAKQfNF
SCwxf76sqrXNLW9nUY83MsZAu7eBUrXeZUfznIYXsCiyNip4ATfCoHa0HQTOLYUcXq4KfAhbCcw9
aSlUekQ0AAJX0xv69BL8LBeYQmwvdlGEcmveUxbhrhFlQZ3hdiisLH2GfQmxUxFxYMu8LyR5G/oT
RDE5NDIXuG++wTsyc0tWweLBJgydLDqcEv2Siuk5BmNCm/IH85zXh7rJQxvPb4k//EJDvBx9DdeA
KtWXPtiG5GgkBnmma/w1CG3g2EW4PU3CwiGj4ErjRdyzVWua9b8ZirMj+heZkL5TlmlrTkpMxexv
xIy82soBjWAwGqM/bdHHKGjXSaguLtINiJ2Qzindq/z/2t9EJXNzDbglKpDtqNMXGBZ+pjN3614M
x5revrLHetQ+aQTNGTYuULtd9eRoGjS27z+L46Lv1oXNrTlMY+1bKy8fWs8EXOBzC3a85yzCrTya
P63kLNDiQFM35DmwWqN2ri2OTnH8mK0lf40M/NnMj5UKMzOcprXssfNMz5SCR3tDLSxKXOOt9oqN
1D/tDqidlXcKYqW+M1pkYjGam8WMBgK4VKI6N6sQFN9wFwkwvIalO7n+Q2orOybJnUvNVMcDNcRc
9cFmplh9+pCJDn03cwPwEoQC5Vwk+Ir76dGXOoMOkBCWutsq+ZJHfQAJtvBADZA8fIefwwHbkMD+
CVRwCm3/B6JIRIwQWk0ZfjRINJ/DfxWG1ZThRcXOGMDs1l/qy9vH7fbbMo7px9JY7Ey/v6xRWzmL
YKtLadiPbSNI1DEtPeyEWxvQFKJ+t5/s8JhJIUsf25k+vnfRpS5u8xJej9sNPgGABaCwK9cDC2cW
93TXhZxlJfju6fmB2YT5FWo35OVYJ8mMnoAFMZ7ZIum4A9jkzGSFby9x+buJ5f2meSQr/T9BZ77x
2MLgClGec0k9g3+MyF/p48SMr+07SsruXJRaV13x4vAaCB3+w3jWkn9Gww/BjCk9HRqJfqHb0OlD
Fc8NdDEITITI4JKNTcTamtVAzs0bE1iBHZ9YhyFur4r1NByg/u91Aetd6lJukI1DWJ50NfQPbdRs
YP2SI4PgrOJzQLoQIvr98no1+TOcqradzHL1ClWJSjKZR8y72auWAvomsVETkN2UkhDI08MnV1Eg
CemOtajDp8n1EHbZnF/rqxoXrFuicAjHIo9VA1n6qXfEZwwX8Xs7TniEEidMX1Sfrk6IF9goB4qZ
uKC27uoCgwCP2Eqpg7yZ852VAACbv9GXzUqW9EJC9m7n7q8qRzFkVGdfaETA4KJl40MW0UAKkaAV
KpcR0Ce9iLtUMJqCbgsmUIjMjutum8zHIWHguYm1SZlI2zmsNOm8AKzIot+A5QCu5zYIVsDjQpHx
wdEB9QTcQPAboNg8TcokrtpVZhAaKcPZoRxV+l00X2vI3MpZpD2ru4tO0MxCJ6nMlD1bCxT9vnbz
jYAn5Z75hmJyNUZdJofsoIs6XfVHrzTULyqUoU78ns0Tqv/SmfXgE2JRpNLsAHyUUdCQkc358yg+
vskLfL2Wji3yteU3X1tBlTTtki/aPIDUUZycCNSeFxgfUYbRaGDpDTMYecZUZ3xx/afnyXbImgxj
0KFESAoWY19o+jCW+rFP1s6c+pGIOnf7sAnY5UpE1L/kJyuKPJlu7oEo8bS1OC0pM61TfSsxyXTt
RlY0rY3IaRCiK3Yd/8lJ3Jt2f0DjEmn+Gsi0V9kWxzP52MrLRU/+GXGcXi2/Ou4+sYagzWfIdEa1
KlcM9qestlmUZ/G2K+WpjTt8Q8meDMIhANlkMHzaMMR8q54JU2Q/1Bo8aoZlRsvl8MMHWeo1gxUD
T3FtMePRk9lvAaWDCej+RO79HeBx68+gmVGTgo9j8lYBgsHRaS5yXC2n3q5ruF9dy06oTPQKO5hm
fzpB41fhzydQKH12gZ8PTavAt1etFQNGbrQdJaS1Bkd1oz2YHhY6zuFLzJxn0TbFm+Fp6dPG7xkb
eAhQz+n7frqH4KhJDRY0isB5gxJmRm3H0DUlOGPTvNqVN1pk2d7U0SMH0ptaPUt7IIwisSkoskg9
l36ZQi1/Y4+sonDamkfNV+qNR/3HIhwIbR9bhTOBZu0uDRF12P9/4eC6Q6SNxa+uWjkYLGEw1bJT
cDFsrJww/xOsXOlhGQqYJmUk2x4x6Z+8xVfT460G29K4WhMR8SMhXIKI3NdZ7rP2ucQkY8k8eSb6
vXSAK9UKnsdVr0zTWzBpJS861fnyiaG+xZdX+MlIzGNFiBsw4DWJXWpZdnwh9nUHBEW58jskgY/0
cSVUuBgxbuT9umj6d6dQa9vn89mu0GlD6DUIvPS2xfHM8PzzhtYi9yp0dDUGiSfzr1+An4n2tnq2
00R77apeNSerhWUWYnRmCD5cuaKpxyfpgaEHDPP878k0hOGUUcni1d/Uy5Ub1n1mOSPb2i4zVyv3
XyHe0M0qVHxEy0Pon531kb3DMv9oo7DNDnnkN6CsGW7nYdcmYfzMPrYI/+y4nNY+4frhPpkdlS0m
jqXJT6RxDj0Lc8ohSLtBz2a+ahjPhwmtcH3isr3lgLH2VGKhotw3H9QpLQ1pH6+4M/iRSqSWPT6I
Ok4roTPwP9YkbRnqgV55Z0WFYpfCD0lVzs0WJP4p/8A7NkTxhK2pB/4CKA6K9fph7j3TFrzaXimS
kTZPHryHBE0BOVkAypVnSs9pteg0q5ZGDRgE1Vy5FtmyA+rm7zPzszz87+hsM316FAdukPEukiQQ
KDYA8mj8pQikIeFUNLjJAkGoqslU6SyBb+gd/nMUlkGCBNhTIkufCEL0bSbcenGyq1vbpWJF9kTO
BvrmIPV/e1fAxQhol1d6vFS9IPZhJx0SMq9gLbTyPRjqHDKbcj0TBr8sYh9FGLv23/DViJopMLul
FRaRSMah4yN+PxTk8Bg8XoSlpG0QVjuxiQLcLe2EzFYoTc9ab3d2brZd5y2QFN0TqXQg5LzkF6hN
mxENuLPbMuryHjn1HtrjzGl1iiq2h1DVKQIq/6UuR6/YMgKbcEkueJ6xepQ9HVZMJcWNR03lZ9L7
utpsu3POsuw3cIFZJ3+4guWXs2kdYbUcacjjSAdraFmPA6F6KVYv357Op2d/gsIdrdI6MP5C2HTb
A71SuQjFj7ORVT3U85VwdWqaPHVZonGn1AhXnGQaRRkxlRFW1J+Smh7/RHUjncVdN0M1S/yilkh8
5hcVvHz2GRNqb0JWaNJD2Td+b3M4VKpbw1+LHmlbNSAkW/GcbjrBcKx7Uf7XQMo2HjbNVvC+yXdO
H69vBQ9eha662gimKDS96brQwIpnwt6wvnAXa1OA8cq1y7Cvyhtsl3BfuRz3/1QJjhhNKvIZFhKA
Sa9E50uy2CKQRaXSbzpIrlyzcGS20xGTPdPEgjKQtLJXy5IleA3Ifmw2JtxwEApQhEErp0bm9phS
/sT5W8qtCQhIPS7jIlN/k5rj3Ff54gcTEjQi7NhAdPpTARZ5sxL+j07InhGYn1OFqyJ+0uLnsz+A
5PuGnR4zcI5FhXB8msWNdvOv9iDoQujuUOvFn52lJ8drv2sRPyvDQcdGq7OIGs3eA0hZSGoBQ5VO
jWHojif8JhR47/wrSKGuKHbLgBzad7u51InyCWw9i9RrUNj8YJQaz/EWbuAoz8TiAjA1A7irPKI+
z3gHwz23iQx4eg/lqQolN5NB1eWIb3Ysv157oVALW3NoHZKUdFTxJF0OMHteCdci9BYX6dUOuIln
GkIX7l27ldXknRmZ16O6iEgU9moo4ny6mK2RbmkJ8rtLPX4+LFSMMlBklfUluNeEdKR4Su8VJrlR
22vs85VqjyDvAuelcovKxQcnsaFlXl6DtF9c3vCamXi3E0if1EW9AX61QPOItDC7VfJlOZKTuYCJ
kpywjYNPcLdPyWM1M/YZYVstdZkDdnI4ymJysxe8en5gLrrVjgbKZ7bkzO/4WkZtheUfhrjNpy5L
JZCiYPjfiifvYzXbkfbOOzA0u7P1qFAeCChGbwiIKDtHysFLhECwmzm9ElFkZJ9QsjlkdTi13cqd
goLAdoGnkz6AUGaIB9xG8uK54uaC4TkeUBR4RlAUTdioY5/abDFmUx2NFAB05rVW6OtblFad0Mc0
ehVaJpYMWMVk36pBH7Sj1J/rBAQVQ2hc9BjN4maD7XAnTC9g0OEjs13ITXvF7UFqXczdALNWW3PV
tUM+TTb1PZL5dfBOk5Ipc3FwSdhExHgaMdsNCKjxhog9fm794+3bvjnEsZz4BJtBoyZOsdbGixdH
c+zXEHuwbXYV+dzosLqCp2zOd238cAT5Bow3DwbozPl4c74551p7T209tiOjr+PomgiGYJvgBX07
QCD7OYOpiMo2paqfeZCwVOjjp8j0O5c2UJlTVDhD5XlCZs5LXxaEdTtEAxNgejkZMN1OpU9l3i3V
px9Ik7a8Gix84FuzXu1g1eIgmGM1d3AhfEZKOE1OSWsqkI6SufISGNsT06h/QZ5+KCdoGvxhrBYg
MyB0y1ItaQ4ftIeVICC+h1vbU6TKUja4o76lqSSwg/0UH7v9mc6ttPNUk/hV8vwxO7Cfxhj/sOS+
b0S2B6NswnR6hcKJQRDWgXIcchQnKQ7mSowNg2LbKAKPm98+gDGV4bq4oEBoEF4saXVHIrL7nsgr
/Gt6EeblhKjodMG/FZ0KZAfPW6GHmKoUzV4cPueNLxbjsA2klEBFDRdsmcYocDMIOJ8qew164XtU
UoITAk7iKggsRbOHiKISNNCJYeBP7vrGKaupWuj3j6s1rLfLZ5g9nDMuMk460vOjEI8fUi7rRD6J
Zl1kfOQyohdnJ7LBIBmEm4t8NOPS57sfz+3tS063K9c21A7mwlt2JZVYo0TvID9nVEKQHIJg/lGY
gMauPyAsPGWkPgbxzNgP2HD+3wKhV9a6+mLqPX5WCMdiGPN2e8L2zXqEYgHRGCsLXNikr6U6ck4p
+uN7Uw4valsNb/Y+VXZQupCh32RirQGKxf/W1VpcuhLaKlxaETwYvDImi2xkut3WzS69I/G6CCmf
D73B/lEzPcZEM5dYIlgqohYQLmKJcEBryXxo8j5pdtVsBOyJmufTwPku8aaqE9fy8NEVDzYSHfHS
hajqUs31M/kt82P7Uga/PmdlI4RH4RSBGt4m0RLnjmaGMbVd72LaKqfDiTmy6FrmIHM7taPSG6yR
Jz1ehUG/BNvILD7ax6XGPImRzRFpZbkpTGYfuhR1K/BV/SUO+7uBuYYSUE95vDNrR5bUifQVMNsP
zdWUHe3e0v/8SACcZbqx+0SuUYsqvuNlve+nrgQ4KK6oeCR2IqzJ2PoRrhYGkIXaxGT8u88SE5uj
J1qKQXqoJM8zLGDYZf2LK9P8BKPGduVHjCJDoPxFI68/3isME6sFkmmybv5iL4Ne8nDqpo+OCzz/
m1bCwQGnC0S0ibpk+dQbQMBCByeXHjXEHASHyzdKbvqVHeseb+V85wZAfuF4BZrgEp/2byIh/btj
6Eq+Qib7We5+zVWIA5DKJHWBfkl03nLA0ZplZUiTiuf+lPfb95p95YeDrxHriOmSbC6c1e0IFAwD
2g99ZapDw0E1BBOEZ/3GR7mQ91Y1gWcPJ6w0g1pBmR1pLTLeE0xW77G+h3P74Ma5FIF9cfqxlrdG
esTZAsxN1u/Us+o9O0OERBzOf1yBH4eOEoH7Mw9ihIfqRzqE78KBueC1AS3U72hhip4C915dNjB6
Q1UODjpf+PqH9HD6pFQaYCiZYe0cqD1lSRT+5AvlSOGYax2pwHoqi1h8WraLleZGtNc7YqGSEgOq
QNtjROJ4G9bLDtWISxwByIjUYxUfan82JZgbrbstCgfWdFnQvqhJ+dwXTFFq5ePT7xKT7PrQk+6w
UPVgHz24stxpT6x2LUnsu7W6XyULexeQhwoFlg/7kVie4RzcboPiCTcy3X++vQKO29n0kn8mLUGR
ZiNi4iKBvNO/c5nVL9U6FAWBijeFQGcHoajGszHs5QZv6fN0MDlpF3nuEkATILFK0x3sLlHK99X1
Fr1NS9G398yuRogAki5PVkfv0AWjWt1AePQbLN9WzZbtdtWRDBShSYb0cLu32nENx/TFwaz8Koxl
x1Wu/RU3hquwt7tpCuJFulKbTsIZ6He4QLsoqT4DluQlupzxRIC/7NbyKyqOsMGzgCukVBIU03H2
CXroa3gIpzia7t3p8zOaEH13Bc/q3NP8sZN0PDcQE6pZJmx9VoH/UWhH5hKmPgVOii9iPjU2zMaJ
vSOlppbfnP/T7uTKxk1N5QneImIhTi4z9EuMLD5r3cQen0Wol0Ky3PV7NjOq2vyjN/1pMQsMnvH9
4id0zS6RAGzkIfNzbILLZJZIsL1/pT7kkB8/QB8IIGphnESD4nwE81Ui74RfGNaqXhRFeoxGrNRH
4O3W8jQ81RtinHy+GUZYucWfFKX6PjtkCFUYktqUGc/L98APMGtIc9bITWkf+10KJEqrl+kUwf6j
pCUnWhhZu+jZ5+Ww8M050ZL4Rp4xK7eREbCMNkzCs3f+XDkiqItyYZLojXeiVj+9vEb95bUeqK1D
aANfkfjk1gNLrDb1/HaHvCHL935NGyBoO/MFDyfR/7nVrge3fNTU1P+C954zI5jBwmmmFSpoWymW
YVoKD8hlQXzUbYr4WlPbDCvcfv6x93GhDNZDMGNkxnFm7kngN/6MrOSVJ/k7qsW2ddroZH8bBIiw
w2pbJRZVzUozRNbwwsnc27pRtOicETF4ID4gkQJgFJgUi0oOxWoXn0uiB3XfRdt/Uc67X9eNTTZ7
FwzkIj6g68fakzlnj5iIzu73RP6y5b8CrN1eRbBNATN/5hQRrNBB9OXupcVGqDzZVI6uE93YqlU+
Yl89CjdpBgnTPXvS4qNlJIVftzjkZcDr8AtGEQEKk/jq3gSaB09EMsjp42LYX6AD8ugxICYMo7eh
xCYKSQFhTNQech/KIihHIb4RoRdtbL4cw9/JyWelm6jPPTtyvWTHhVHXijSniwYtPON8+cr1ESPJ
bZiHTGIPgZAblsGUkPzmakLkF3F99DlABRF4MAzk3smMINgc+q1pUgYs68LN3pJEq+k5vkRyj0l4
MQL99v92RhWecEtN3mYBXCCHkNQzqE4K1eVAlFtS2nYkaJ4l56IwsL75aOcAiln+NE/wTTIjL5bT
0d6g8lgzs7R92ZnC8pq9J1kiyDPjyXGZSMm0z14oGA4gQR2mgbTIQrtQCctLqnibIbDdn2l7KNGj
zcjFgedzXhR6cdlQgXH9xbv4SITYkFF430nQ6v3MKLQA/2lyiHNFov3Vpxep7b8IhRL+AMEsDUAE
96mpb9tpfGE4/uj1AxEAKo4kM6ynm1O7m6iuDprXoQpmP0v5Lo5gLXlm2nNR2GsolkNP0GhcKtm3
bjweFqCPDbcpP1nRXdGbC8oiLA86fTpTAEPtc3AwDHktqKEEcOlCPwf8zBYKKtnFVRqspvp8K96k
2Ba8gvpY4J7LMsOg9uoiq24VoN7dH19pRSNrojIY48r4J7JT8c7CcUK5JkBdXuQeyWYp9LceWpty
3u6AxZBpy13qnLb8+o7TB71rAfWXzivrlBUZaZfUN69g/NaMERCcpWn0I7+BG0h//4dtfe9N0okM
N+m8GbAVrENWB1wHq5BdgOSdERkP0WFIn3fckmokbhceFBbDH9X1rf6SdgK6URUVuBmvY6ZGbMcH
l68nhYi3OoF3kcpXuHmyNvD48ImsJC9hUvmfE06Dv9RS1td1TbBri7AVgMsXq1R0I/K4/1I4oc26
Thb2kZM2IZlzahQFKjyFG9k7RrS569+FrMXXhPqZRTsIbuB+w93x0bZmrooBFSvyeCfit1GwElYP
P8ophBgDO36Pxd4cysgJsf92/jixCnH4IMDJBkOeCym5sGW33uoLzNh6IZjEU7lTDyi4UZ9a/TEx
eLAm0d1ZALSx/mW46Xacdd+FimF/BJNOxe4Y1SliAFWXRVUw9pthoB+RJrL7RdGDcUM1YEZ0mBKX
bzpvDd8Tk3idj1NRd71woIKjhEQluDmS8vLP+9BX86ekY4gHGhgXb2vE/e44/zc5Amu1MuQpqei6
16SjH05pnWqzoRSpF3lMCBH7P83f/z4Yhw84yp98qTCIcDAXW4tZdEULMG1yIyqZs+42rlFuFHg6
jhPVzxllQV6A+IfhQAKa8rA/RurZ7+xtYBxIiBRBM6jyU0DSK07dnZU2LEuP/G4yg8TQOPL33YXl
5BYSMDRfSWIOkM3Cpwhlnr8Dvb3e3vrCh6+oeta+un6QWsG9YCIoJLaiHmLq/LdgINov+NJpuhhM
3nnpy2h0X2TG5uIhG02DZYMPHYPcM5Rhpta5X9F+IHzdduzdCw7IJu+oyUhElWhVx6Ze8AVj0EPP
//93TJ+CGYkFCLLjtLwwYPMUQ/kBGQHGBB2AQzm+vc217CHr6rzz9f6fBzqCDDUkm3ScwFyAe8CP
QEkfL4cq+MefpiRaE2f9Qe3PB7kPD+rTWGirVIuPTZckjJJZ/1N/OAdda4H1yLpzD+hHSb6NNa0M
pTJP/U2I2kmvPUHE9Z9Dqi8vL36MorfLXAbCyBd4rXCjmb7nOlqF8zPVVvUAn6ClgRx8eAcR9Qb1
9i0pobwve70NRLEaUNzjF0kGqNfhDG12WJX7/QX3Ihi0R1l62Mw/mEygfOrPSVbN9jX/Kbmtio8p
en2rga+fHOuZhdKMQOPgCEFHKQFHNCYzQ0PixllR1+jox3xFVTVWw/ob+5M2nRE9hdr36gRgTOda
znnuFOwvcJTsLCEjMWFPQJTt/oZFrYjE2xSbdfi3IH0iQpjk3MrHYhmQVQ7wV+6pYxC4Tz5Jy6nF
IlCcm7BsheUZYJD/Z7Vz6v7EuvE7/He6gD/nmUosFx04NYM2AvX2FiC/jAyHaO/x6EiWkDnhdbQS
VjZTOahcaRqY7Qny/RnM4C+u27+Va7mBMpmv9KpuUd//dw0Nc+syQCRD7n4T5qMU+9rDjbJemfi5
qVBQ+2FtaQ4NoBZPB876qHF0kZtsqrnroGXC7ghaGETvyv4CCzMmmw5NBBaTBxyq7zQZ3JuFgm6+
0x7h7Qwu4QW6F/OgOJ9s3dJprEgs9dECGuJDUx8WFI0RcmzFoL0ZNJL/pciAv/jjsDcqaUEvyPhY
a5y2j4XszQghzsj4Cwh4XhpeXjDmk2Th/Bqe0Y44Sl0f01zGHz5ZZ/jfKlayK+r7fV3gXoPxD8Eb
4qtkaQfP2XrbTGZJiGdCJUsgW0inQFzM9xalp/cjzKryrFY0/2ZUDKvzjgAbf6ocoX+Aot3HsHnl
t8IfoIJ/+LcdRtPQRGdZ0980JQ8ehdqpYZRJxgcFOhaGCl8T3uA3KLhC6UgJMrzO96N7isRLqgyN
E08JyrtTfSXt0hdiGrFlGocaJD85tMLtssPrxKE6G/SWNitWHGjwNwT0SWzdsEuTQYSLC3yjPfj/
d1WcyP5Dpxo+irusbMCyUu8xekN7tYaz8WqJjtr4rysvwz5EzH5mV5mSi5Kv/0QRnqFMMVJCq1S1
YzeE2oPRJrwoLC/J8MNzRPazA2e3hIf+wrZIfzTpB6acpP31KbD2BbDTVXOq7QerO8rrXqrQqd+5
XkORotijFxq5Ra4ZFbm39g99AXWCg65ed1Gc8f4WU4mP7f9BnYgbWV7oURVZ+eYNr6oIOx6Gix2B
ZTgg5jAe94LDIdtAh3KzcHilAXEa2ewzXGCrtmmB8E/Nwf4hME0PGm6NCwdu0Hbnq68V/TtzdVXK
ZQue1Ys1S6kf42LZ/8kw4BjuddDod3jmSPiWC2/qu4ca7vrrpZY9iNWP2E3OB965A8FJIDp6DpQe
TW8eFIX02ZCInnTcV258hz6fGrZ7gizD4O/WwVEx8ujQK+qHc5DqQmsYlWyeYugmXHhb7+zQJ+h+
CzzadrtiixII9TaqDevay1TUwD2b2HVG7qUiTzPaBJ01wlpkQ3sbLCQ/Lt7y3CtwRowdwbnXBmBb
0cYQedNXDhJ/+wVcbc/HJf0wBWl+6MpBpwFN4uM4uxwztnVb9rTaOgB0btUdh9Ol+e6zShrO1ELG
AdRaztT2YmTGEHa1wWrM/A6RvuseERCGaDLT9VqKxJCi6D0Fk+d5TBchfLUOCCnW+sBYRFxFdMhj
7OWFLG7t6lC7XtqbKtEhFV2y/ebXJSh5t9aBME65GldBThwec3uzXupxia4uhqYpK6URqEj2pC5x
2lyrSkMM3/46RX+cT1jSPdaF/viENSKiIZifgkE3HwHyT3aMReTlxD1SQuKWdBCz84RumX/v46tW
mxEI9OFiHxDWTSjKt0fjR3x5RxhiQqfZnRSbjNhlcyKjTOCQsEymKhpkU8tpQO45reLNjosonK3a
38GoS2D4gG3kgW2nISqvmToPgLDZu+cjpQlXFPFTh8hYzTOX8WWKHruP6Z1RDkEPW7lneZzvjEQr
1Upnq0Pz/CI8WwdmNm7pV5KsqXFp8Z+we8XQmwdQZVjsurofGACftXMD6HDLbdc/A6aeTNe567r1
ikp/xyHkR5vRw+fXVRmxdcUWY8Or+7UgI9M7AmpsURG/hKZCHUUjUwShYJjNNB6E+5fcpkBFvPl1
eXpaPacR4LdX4TFdq07cos+9NvokHCb+Bb8OaAv+OHHC4Y7OZRLrJRP5okPjnTN9f7LnHIq17cRj
mq3w9QwZQLVaoDs3aTbuv0621La85wHmhS4b7htLOPxNoIibd4sEjuhiMsPyK1ZoqJp9gnRXuLq3
rJY4YalLlB9fGAHahKPW4aVs3GF4Por6hpSPio6Y9eM99GqmLRSDBZ3yWXEE1xy/2sRM8yOnGQk2
jedgoP+DLiF+kE7PLx1CTZuDB9GpqOfXB8qKLPh6Mcw8np0lkTEQF+4ccgRpCMvgJIbXGJfcJUKM
SnSXHtT4o7c1FyoiqHiIAfoowqUSgf15ulwYw0Jly2covnjFsa1TBB47z52q0LTxhxaFwk6H0YeR
xoJb8GSNThrp0G46RUwOx8+lUBUu18r0JKYewsgaZzJknr5BAR+yYtJADbbGDPy8rxP8Cn1UDgs9
INCjGwqy5XvT8aPgx5Tkr8IpmmDykpipeJ2O1NV6K+VnF3P/Eb18192pdKm2i8H6IFQKm76JDbXO
RfoSNflKYKTWyQWIbYi330hx3TQ8lE1NlSCy64KU43suzRJb6nRIPGEZt7U0pnpPgtu6YsmPm6W/
tXdrlQRkDKErPYeDX7jlaWQ0NzFmHARGvrKZHyn+yQnxY2W9WHpIyVf2O1Z5uu94p3Bi9mJhSwTy
e3LptI8RQbOEeKGBxoVM4fIIr76OxE+eS7W7Yuu16fNDIhTUcICtrjFaHIDKw7AQISW7J40zEhgl
bgVL4sD3rWGAvs3t23OvQjaFkJPQoYx9gKqCbRQBmNb47+35QOsPFf7Fgn74oNOGr3Iq8gETAzea
ViQqvX5SIEwpZdXPmptW+bhpW2/7uykpk9hQX3R67a8h9EGTf6YhRQ39pNREZWKGcT+wisin3IDb
Lqa82h8AYXMTUTtJiFTqC0oia3Qali4MisfHze1aDaBuket/VACejMwBARuzepWJzeHC2Cbwt2Wy
JLytPLMjky9xS5fagqh8DMD4My7uSFsXYlUYCbRIwViLz3OzJw1ajOeIfIbYVptLyIg9XTUiA32j
ywr9nHRLI26U9ohW/KaJY3PBKjI4Wd7CqPKLQ2TJDXFBEjc1Ykl+ybI8qe4JiwO1ynUYRKGCUMKW
KJhhRBPwIG4Gh/R1KgpoE5M65IHRmoYx3lGhgasFBQUBHZxE+Sz1Hx1zTU/tm2IRZIcEGRf4PyVD
mDN/CJvqLImHsMTMAqR21a+TeqWznKZhayfNd008CoCNenFB3L0ORI914maowJgw8NzSB8yE2BZ+
pFnsGuDJL4uB4328PpMl1tnzaVHMTFunSpTkWqA4fOVPXNqc5QOwxwAKEqCfowcY073/tYyw0+zg
q3HKJ/1UXfV65RQ6YgYu5VYI1doW57RPw6BSVpxGG1UXEPsIRFCSUXQmCaVY23q4n9xc0CP391nC
ELIOmF7vvtlXuWSLDtCAQ1w+uBpVIV4sWGmYqH07LRa5mlrq2PvdMoBjkt9sPKxUsOFcHVIVnz1T
iObL34c+Wj8pEgN/q6+nf03sZBkd8FcZAR4/kotiKNNOYSHDxNjuekS5ZtbMpKnPm9z/il5iSyml
BTyBuH4mXLHiuJwOmU8xBWg4nEexsy/f/D4BFH8HHi9Md9obXDd9dWyl7vqLLB+u/cYnnbKe121H
TYmWD3AW+MaFfnOc7VKyxRM6Lfj/J4qZYCWnnYrYJfC7kTC2r1ZTOZuD45L8DYnuwP3c8+x4up7R
aLD2Nak2/y5hUqkfHz+8+59XurVAp0DSfy7eLlAqp0OdbDVSOtcCflobNw7QgXtgxWFvWqrtmJIK
5/Ccmvf0WoV9LY+VohaQNqHGc02PDsnSVtrl6GSkL9fsdw+i2HJTsduckmQ5fb4TcmhbLX0kJ8j4
E2GrHhxEv5rBe6Krf2nQpgdSUY8Xuv5usbuxjnZh8Yrxuz67FiB9oMUENZrmCAuTNa9Kj6y5TuWs
A7bOu751D5rjHwz5qi710Vc9bURjIcvCdJcJTNr1Id0cZodCQcRLRDlR7hnH/m2zkTXxOWNN2XRh
UF4btlzSZblzJ5FoklaytqRf33srkwPtncJLZdHgkPzex5S8OLBZEDFBzFPchLIzVYXwxFEZYNqW
J8QfIqirtKs6quaoQ2RHXMyWy9HyjgmZU/hWeEH6aLnwhDFrgDTSElkLeRz2SzrreAqC7m/n5XYj
STycrJJ8jBRvHmNMR7Lhbfl5bJgVFvZL5i3SqrCTOIxxOCZEM2eRzyFkqZi065xgr5RazNla/Rg3
jlRJ92WvbP0NwVRi5K/C7GqAGe7tW5Pa0Lt47KDSCi6JFT9jjeQEIuYy/TLtZYbnvVL5kvT/oFJS
yO+CTdVW9k31+Qs5CZoM3/JaQ/G0OSGBEg0naFkAy/axrp/5H/uiUpkrcn86KOiS1xtVS7TwhK6O
rNq7HPj7XXSNGcxfQrG4Q0gMVLzd/TioHjaI3QWVq2ytuO7X2vznlCf3mfL6TNsJhnPl2sZBKoBk
t872juI6NcrRm6lKpbF7lORgGW6QvCOQuhwSKjVZcqtoBKueesyf443EX1THc5+hWw1VR2/50Due
ameZ8C44YKlQ9gRXPcVMZrrv3Ako1i9+2uYJRBwleucnQ0BJuCYNFv0v9AWwynDPngeOJmQLOqai
TM+NHkeSEqFAnfR97J/hu0LbA+lpK4gSeQEfMNO5c00MRQs/gbKcJS/veX6KaG1gM9PzYiGfOPqd
3huRHzdCK+T4ITcDmkhdpx7bOXcMwgDmXT6WgtArm1/QlTlAmnKN2ty4DU70dzDwiS263n6Gr10E
F1Uq7sUn3VgPuv0NcZwPT3yUqxWPsso7UF8O03fgGDzW4MnKef3qJjDg1K60obmQj29AphAT9Jrr
Cy6MhXdQt8vvsmrH0w0BI+EWoArVDWdAx34DBy/yQ4BMRQP/RoQftCDmxYtiJylR5zrjLVhNQqEW
3qYPtN5d+8jzBrTivudYZCc1np57kxJhHaiv3uk5ELTUcTUM38ebneASQMbNfR7cWqyPTiQ6YKXd
cZMDde5tYBKm9cW3nrai2N1+5fTYAA7p6YG6oeymBjn2LJ31cU/HfgZsAX2EX1tPfGhWDlZKyj0Y
PJ1Z9KR9ULseqnEFzAeGOsj7oWgc0u/1RptU512hXG2Wdwa9p2LEBJwn4BWpAgKJdDgf1jq57zs3
HR9nAtWxUZpvCNt1ii51+2ImLa6ooWRaV4MhSGPFdn665pYOdQRdyXP2VgEX8pMdx2I8lq9/q+VV
LMNc3zrpKKxk63e1W0DcvgIf8epPk8egqzn0q0JZlQW64IGOXNE6M4aRqDimWJlnLvJps8Uaowam
3VJXQjiknW9zGYLTXBAVBjOKpUumwnlTy1WbUnnHfBc+qxx2gdhud0/cD+KvWOQitRC444s7ppy8
pMDRD5vfd9gCdmen4nyeSlDqsIeok4323V9i23U6bqebZ+UPupHr/YGYT8YZy6fttUHJZvEbLZOj
4Ns1TuZ35KD/Pfco8YXjP3xguYUmNh2tCDQwAWZxx2tM4lcCSPm5oaFAXXunE7AvjPW0F0zcXLW+
x+gzptK6Up/JjYhwpoEFtavnbhdMoAwrh5vyleu8CWMg/Kb94IfDVsPvi6K/j8a7HVI0RW6uDiDl
1satILxaA87tBBqBzVxktz76Skuur8qJakJnQ4nooarKCSXsXGoT0sTC5gb7QUuOoEE98i/RWIrL
E2kWU5PPG6WGUjFF3x2i4CCk8loz/O1wkKkUmAZ+fA6lDCU/sARrOka+LpOPiXLnx1DapU2SrlmF
OIkDj+Z8dYgQgshDDT9FCImvLM1tBOEl3cO3h1c5Iv3IgMyoqV8/Dho+SgCzOXewUygRbbKG5wRw
vjBTSqQwrGZ9VF3m6Zxg7/JFAxL/LGeQ1hlleI0P9Yy1NFpa1EhqhQu52l+CBoWT0RQcfSvUgmOm
tisQx2LOKOrInO3wpv7ioJ+rWpETTJEnbWEsLoycMtRwMizI3gm2Wo/imD1AuODQH7tl4PFMkzys
2gpoibDBXQQtBTNn/EPl8AXAXmv/5oYSqT2c34tMdT4nZAhywKAaxgJNq90eaDeedXQq+NBJjPMp
nPcXdqYuMp+33BkSixxmNqwyStmavG2ayqD/w8rMsBcAG04OR5lr0b7nVhGnsFEgxBUmgbQenKmo
KwpPb8qcmWLCCQW9ip8ltUhhGen+tm/AwxAU5AtjfwQ6CQ6XSRGQvxA4b+VBrZTsOp4YDI0xTKE5
BeWLIR1Q4VkBHOMc6UX86Lr+B4OWmtnxZBqk/xzEApYtQQ/MB7uTjzD5Nmb+y1w1x8QOTQIoT60h
Pl6T9Ozpy6YL3Ry9w/r3lmoFPH1EhfXvB/A/JL+W6bRUNKwT3oAcUNE9yeck8YawiDj7NrZj49i0
pBAx6IzhV2SS3ck8lSxrKMKKqZTpGa7umDpoRsYUIHwcOCAUutDPxYwlmJqIxeLh9kf3f7w/FRWJ
COm+zOWIcgdaej1SsXX66rR8EB3kFV3QmZjXVYsfmrZbIpN7LVOwjyzM7+sPFOiRybmU3YtnPC8X
omahg1yjUgM/P5jgV/9jZhokrGYrHl2z38tyW4vJaDymPGAQXP5/+bbczFkwgyfB8SihGvmxzLD+
rqnT6m8XIneHmXpuwvUA16N+mN4W0aXD/GGb667Cq8VhdhHosHOhu9TVMn7vPlNgkLFyEiuq8geI
hrSUtRm67E8ks7KtuqM8vruhwHrzwd7esF7bBRYUzxeqVl+WClh+5PHLNR5/oEobxE/1o2KTSX/s
/n/i5VFrno7iKGOC3CtUB5YEeEcaHymx2b7oovtjYxlXklLbdebOykrJEBCsVDlTikR/K+6nsk8j
0RaVyyDN4q1Q04b/ynV1wcyNG2YmPxwlLEAIf08bLL4wLGBxsZUkG4dURZgt6GpnZWxh4OUJhBYD
d1w13fEre3Gejwg3AgghIWnDb0cnAmFgY2lQf7rDEhQ7Qdat9VhVD8fk+RFnolrgIYIpxkgeia/2
9WiIzLuDiBGk6NSXyz2k3DA/XT7SKSAZzHvSGe5whY8i6L2feaVR/aSxNArtCf2MHpWaO6pawoti
GK9YAkc1Hxz0k99wJ71caP1Ok5iTk604k+i8EHbAQefhytOrlfYWapYIxBoLatPy7f3dOQM3pxEf
Wf55wCfQOSQtTUdN6TGeJrZlhWfoHOFypZdFUzYd+nNpLMNH3ory6d/hbmPXhXEAJGlOYm8zvKBb
uBaOvzN9NHsRK+KAKsej1iwR6XOcuUQeQkTjnyUrQ2K7Gh8fmKFjzsC78Qy12xOQPiOqMq7UGdn7
pQmQVDuI13sukGXSTzV8LO5/x3z9EgnBY5iTUiOlDeU937duM7TgqY05OT9f2OBXHmhpLY2RSuPx
2KjP/aJqnzH7S/28rSZ39saNXXqInF2csgqT6nNW5Ic/LqO4fhscRMc22pQ6XVSx+wbpQzd7ERnB
/siYz3TVBxn4zW1Smp8xrS5wZDywjC22mdSg+f2L+59M/rUoYd3UzfEBoED/mNxp7Bgwp4dSC3Je
WjVnLZYl51meheO+24Ru55dV18ymO2JaKHW7Zji+303Bt4by0Cnmv38y/QrjHaqs2L1EoY3Dc1mr
pPWSt2UVMbkk6X2WbUnV8Ps7G6OD81HXd9Hi0w6tiwJmTwolSs96L21VFlOealzrtKeqK6aOulxP
LCP/WIQ9L3WLn1fEOJ1R4n1MIoGtuUwZnhpMRuh8os2o6TWWNHLodOdz69RcxiZDjLWfvXjqobX7
RtGY8HxuJj1901Nic4bhHt/Y+dBG+ktQJ81I73UHPbnEZBVOG8aQR4BjN+6nbnqXtBClGnJULg6G
LyN68e6snOjOhS/coa3KtGe8EHTmO2ZPj5RpLk7Hpy2MEBVxFBGEG9HTUDAbqFb1P0D2BwX6hkux
q3Hc/S5GutNy6AklZhNbC7stiAYFaAOkgffg3XI1g+KryiiCkD6IrNOheuOPiMOf0XH4h52j6fjN
QpXMFmPfn5avv+BuBFoCkCbePiFp9SQVIUL0hCu6cnP/Bi/givhpLDT7VlAQ4zIAJ5jNf5R5Nwut
08xsDm0+GDZc//s1oRopm5u+cI5gx7VY7WY0iP1tqgjHyfJd+mpFRxGlm5YYoACzM+mca9suMIAE
anQLwbQu+fDw1RKfLIzJCdpJw1+by+bv2VWH8jmYLAJcyOYXWV3WZZCG1gAMmbcYG1DEQJJv7dzQ
P45QshgG8h8HZsSvKiV1kENv+1yiSMU0KOZ2E+8J02C5rpj+Gaz2jQVa16i9T1Vb87lEGqzRIzI3
/vR0pc4YWVJ8rhZi60QEeq4GMGb5+2PsY98FPHZQ9LkuTQaFLienK7G9Udh8yg0i9LLNN5JKzTPo
pv5IdymK2dOtYpPrF+zKS+5aNBWeBU3yudzpCx9gLlr6yIbyP4lpPpbLBfQHpvApfm3BDskvfixU
EDdwwF/GSyOsk4t/qXjCSK+X3zjjw9TOYowOb6OQ/ZnnNvdcqS+eNU8eeicb2v6osxUetnw/OtzX
+FXZwbjWZpCIRyZBatZRSUZVRH538KSAj2iWeNSjBTwunhVYSqApofXKX4EyCfFZsfSH9w39DTa9
7L2fdH2zbupbx92lXyPZHJYxVdkLXoP7IYyK+H5t977yGU+jPoK2Y0GaC/kLfyejdjTqNkHnvBvv
HY60e5sp2Gd29IwZ7laboMO3zsxgyojb8Yj+HGuJcxNKYqui5s5HKcDnJVoc7/6L7pV04PCKqTMb
FToXVapO5QJPQGK0SUrj9V23g1AyZjuyn2JAmJh1nbNBZgVPz+kzCqUsMSaoxuDRHEB92ML4Pwg2
zJqy4lhTlVBMwOl+k4ZwEp1WCVexebaZqfoxB/tg0wgwVgaKILe6Rrzp3tY8J/MZL7CmudyffIaC
inqT8cDGGDowwfEiCqf+PXKR6QR0VmSaXXJ/McBidemnjA2W6mImYp4RBRbqJ2c0HvySltjWwX0g
B8ZKahQJ7gwQQq6LIKYphvJdBGS7RewbjpoXowwSduPHDjB5q+Ey1Hea2PeWmOoxx3rJVUeF8fQ7
5tHtEuUA6V7rEO7446tt+IiWG2xjk0RXHPqkOFnc9Eo9gOas7TL2KJF8mB3/gx4jUPZeV3oTRONs
nGQrf1HuAfLV+bzg+eLV2M2ZZugM1sfNdWAlSQmmYjmvYJQL3En8q7h7DFpeZDPsByUWCGqfl2DF
B0XMhWAPC54gvgi5+M14gwTM//YOt03FtmJzWaRvsL6/OOvEaeJDbrN+RrAdieVPVIPssM6IAOmM
snuY1yAbRllE8QTx90MZpHIh48BRaRjXkK50Wdr+kntvZuzXQ8dt4k5vx8qKOW58PUQXYboGZTTC
IhIqxZuFvqpXfTpBrYHAmjznVPCldEdvFXhNKuAwjLUrFD/MskmpNV5TMCxDx0TWJXPB8WhrD6wu
e8W9UnayExtyMUccxBrGp98UMFAGP8+sOrCYwb0hUf38z2ufYGv0jD86Gj8ocpkROriLgu2/Id+i
erEXcOwxWzEVIBghbbc3g938Gkd2owvWzKIRIrKay0xc1IG8xn5W3RGvWgjkPYXqbi8+9AiQajg1
ix6AMSvNcpgylS/3pu1x1mNGD8QEiCJeoG2jBGAa/qWCttLaO2L/kpjIy58LXENmaqElPGZj0k/e
INKpyAQkI3h0VQyCw5bxN6uUAckIhC9j/j56OYDmDRb1D6CMjrbU75mXZb0c5+frGCkkMV0v/RP1
k0iasm6biPzcyV3X0W+lqxbtENSKdVHZScG6dj1eEl5ECfFhxthHNLz3aQcnjAbbKtIswy+48Bfq
N46Cgmk1UONC/dxzxa3Cd0pGqBU4nWqbzojpyVAq9xg+gmfhngxjsb6tH7DdgUwgUj+mtMuFY0eU
TSsBjSpLHKZApZUklMrlHY+9rifP8TJeZEFfW47ZdvJR/p/LoxzGtoyCYeB7X+MyfHGOw5ODtejv
QOLDyyDWcskBEJoUcPWQp8EAt9MLEZ7Ogo2Jtnd48h8nwcz4qZwv6XM7pYTjJblc5GKSb6zndy0x
VNVrTckLJg/92iZKwQ5lG6SE2dXX0hyBy/W3wdz5Jc0XruPzvkCA0pLtwofltv3s3E0x13bNL5ix
XS7SnmRz7y4LFlsABkKEzJFhfkE5ItJRBak4mpONftGuyHkOMQN6mAsKbulk+an9Hi7u4LQ0YQap
3UW1Gyt2m/IqCT4p4cIK6LNzxyAtnrs34UymPAUbWth4x5z8RXYMSDt7gfQBhzcfIvG1/v6MpK3z
MOryBCutqPt6DMj0aWAvrMJgSDhPSC9FO8z/zgBUDo9qtQ8KzVpcrbKUTDrRy/NmMH5D6lo9LENj
EyqxM+Y8O3hOYpumLy26yVN4oNR6+Z/U+ayFDUrtPs8h4lBfAx5VoDPEOHcbujWdK6FDMKieoqd/
5nlwSxIdxEpubmRxGYDMUNP0D9AsgOXfmmVeAOccXoCUVKpO6lgy51NlYEcM59b9ntjfQL/rvzZW
oNWQRCVwMM3Z1lC/IbSuFTCzNbgb2k7m6Ot4bku+ZNV3WHHV096SEPlv3+MZ4bAEgkzXTtKQjyVD
9dHyGSbeXbeH9E0PXeYymPVzS9xR5xSkjtvj9FJgVgG1syoZuEp7JYNKerYoH7fmD92VfBTXF4tp
P2yMl8KB31V9Td7/OqMWMQrdS+50Sl0JSl8v1xP6Xv+mFUnMUuif7YzOlNtsNLw0r1c0Hzx+o4tB
5Sr3LYRSr/WgBZIoF7t9oE0nkAv3YQNEwY5VL82cuGrg0i1aWzuK9AMpJOMO8QclztocvzcBrVer
2krZqRr466X99M8aviiAYitryCzjz4u99wISZP8mgDCO3OgeaVg9n6yR28V7+mhggd43lCDSS9/0
mwvMnUV+CiinM4UV/ltSlYwIIaPVE8OfEzTDloDYBfUE30H7I2fghO1+b/R2klrfYKbm/PO7+QvU
ma4hUYtdaynS9RCsDOri35Lyapopzkr2CjTCqCZdQ5AIRP42hZe1kJuovg+7uUdrtzvWkGreRfko
69+lrO2P3PoB+cE7daUzuBBWoaSTswkO4uUbyDukV4kThIpn+dlsZCQaK6oMBZk2Mch8EX5p0qcN
sHKjASQ9K9n1nv3xBSjqBXLwUOpGiPb4yz2aZ4bOZcP9Tk1tB+umgBAhZnDFQbxP6aiTrJLFqFyE
OTZ5qYnoCI1rrJwBRVh9eqdsRsAWQk5ICisNyVUcmYmvJbi2vpmVI0WaKxGU/mFvqGuVtc5gURS8
Az5q4Oa/sPZ7cVo3jJKNPh+rG8Bk2hes2F+xK0I/0rygYEWV61v8G68bugoMzz1qOcRdIDN2+s4z
XGcMcmnWfmpSaNsiOKYt7VdElskMBWE7S09HtlKX4MR4CxPrGTNE4LQzx9p1iRByp0J2pfu0zSGR
wqV1O4tKkX46M8oEpC+r4e+JLkYKlmAM9B5RSFuJoni0w0tNJ2xqbe1D9NFErmD94QSkKzDTSSnY
C+11/K0XYYc9JHP35eMpyPlxPnt+ohF2fMahcLMaNC8xBgRjcrj+ayRv+u2grx3d94Ve6Sofxa6z
mEO1QJfL1UXQyJYudEV4Vm+CuEjm+JhCK3h3h8K3x/+AVsWihIiROB2XUZaxYreSlKZMQacynWFD
i9rG+G61g8ilqyozLUii3Oh8lgp9ktBVFKx6PMaTvJh2CbJoOjbBamcyMGCxfF4aoXDJeF80X833
l8zzbypBGxgMbJcMcWXuC7x9TfkQsNGkxR2CK2MoSMS1kN/tSICaTFEi1z1kpZRIncrkOohLV3ui
76m/2G65nMFvbmyMnVHBvVMUFTVhuxZv5mMX51mTKy6Olmmvdw7MMToe5wr7/Y3Ox7xSO4R6JTC4
Y+j+X8lIXCmBoni+wa13IRn2tyP6daVuGIT5q11Y56tEPIFHBtHo8dxVEDEtDyjSlqlORcsICv4x
SlNHMbwzKQFUzZ2ZEjhm6S6VbGMUhGiTBcyqqD2JGWDs6oY9Z4EUbwNq6PoLhijX2k3iNgMU/IHL
XTn2cEnalBxEu6c68IyUe3A3u+ix4NV9In1o96Irwi8UyXQA/oGQPTvuFWnX3sTJX3KAGjAuNah5
PFwES/HMBBuUHTkQT7e7WjlGind3PDdY1RZfz/79chjFdCYQnAybOpMCYxGbL/TiEflz383e9QK8
PIeoQER2o8O9IErtPpnbK+716mRcYn8LZQ4danwgaLooo32pvS/ITG7qvtMeyK3a+rn7TEcGY1xR
b4pyOJm5xxUvv/fWpAOtcfCnum8mYmyYuDDhvKreQ4SG/tivFQC58sXOAaDQmBxOACfD/A2x4kGl
RdrZM3aOfdQqhds8KhXcJD8rb3SNoCYarh3AOUZvWkQDnb0Ze6p8mpy36gHKBadvhcPo2jNkArD9
3qO3NVHDpqxYDn4K13vX2NZKDzP1c6Ae46joumeam4G0KFwu+uthn+JDziUZg6TcJRRc127WfrUR
OoVoFvXQVT2FGLjP0lORUzqHkHyvtmn25KHZG3WxgQyMLxmzkTysbD271TEhtjadaELXMkVbqbuO
RmjSR36wEyvgEHBiavp3P7kjZGambPBF7KvEf2dHaBxMJYm0oRFKo6CEh2ymQBIMNZ87FmXxPgYt
Rk8V2tw/xMgxxKmEpv0sJgdxa9GIlsl+4hYLCmuqOBwW9G5/p1lI0Q2Ciw/fYm8Re9Q0I6nm3MTZ
cCQGIPdXMGQsKm6wqTcM0Qk7jROwg+Tg9FTbt2d4uqE2c/4c148TgHb+KYVEe+aOCx0mxFo1Ubp6
LHcKyTF+8Dm5IP62hQ91D2DiSuZm15aXN9GK5B8/WYB7RaFBbGmCM6n7GE6fmavepgMcaVVXAvr/
RxsrKKQankXunIMCF48jgANtNHYY71u3n6na7jvQxRo4sSE7zXL6lQSVLN5Da56BxMzLqGGPHuEM
19rKuYjbfK87zQfT3lH3zbJzQam3m+g1WrtbWdVuzw8Kao1gLSko0MrKjKs8rLPQJ0QpGjKrcq9j
SBZUuTNMtaMXPzT4YwRPoR9kQqvhXTJSZMz9cwRaOMjEPKI6Qo/4KjN9TXs48wj1H3IAsD6gghMI
qapWkfDGtVVad5XZxjmsooHYyR6QBSPYWVM01r+h3iVVYRGm55lA2PpVIe5Qo2CnEV7uZFx/XezB
3K2YUEFrsGJXCvqWYGJ6vFUsW/viBrudkeOXEGHNUfduJxqR0rBmo5ns0EC83rq92SnbwZ9yX1yt
dSE42XwTMYFozChfvNyl9m9fAhHOrpSWGcQFB8DW8wMGOAkZxd78DhGBddMMH2NiRPMt+a/4uvRK
BHQN9HuWC1b3q6THuGcBv2GOIzo3kBc5fUDVlHFRPIECF+X6qTKfsEDOA3+GkbhX0ac15MCrvrEr
1OGUv6peus4WF1bWontor5tUiceFowozZ7pWEik//xd+oP/s1JZNHvqanFFjt+CHA7uht4kHrk94
enbLkRhEpgygj9lFNoSAhhTKAvuvcXDCLeX/JMqeqg+rS5Jwtn9qDHNGYtSvT/yvwYULbRU6fM6c
xxaVNBoMwnrKHTUe+2v0PXhH/MCv/bDAQlIJX0JtUkhyh4q1VhWqJXRu4NX/5ZzuaV6oIDmfFekV
cWGbfUSscxxz9Wy2N22hOEmBrOPB+/UcVZUU/uZ8gacBJrG5WmtlP9ouIcTsVF2Lkv67aS/Ww+uV
Hm/2Mx9us1yCHyfMpaQHq8RHzrQMKCZCmjYpzgPsXRM7Hyg9fEfzmg1nXhsgnP+mLi00nOjRGzhg
mLWuOu7OOW4OFsQRLx8/69izBGrLEyNy8T26E8wKYJ0DP9qihp4qRScw2p1NmpzlmjLWjRoGBU9F
qAoqTgyu5Uhvj1UPr7DD1sBHAGFsLLeara0a3nDRTuP65zZA9yba90O6SFtsXNk5uZAF7SaVjMi5
n19B3YAxEUbDav+CWaqP0fYxaemgWXdV5KGxkipFnzWJP7/GzqYaOWz5HMl4T+sQJS9vUJslHREI
GYQz4dr5cQNCWyunKQ/NOeYsTpJ7OGNRmyNhDlRuHowaO2lTtd4A0VXBwdv+xgqf2MLmzbAYhjLK
gbg8p7D10c+Hkt7WkwUB2ALq42dKO/2k/aSmGZ/2TybpoCcVQzAR24X4kSHb9LvMimNEvwuH3rbD
+lPQSipJnaxhcCD5kxdMpEt+3uwhj4R5cyMEU/CkZeehb/+Qp0fcSHKeNKP5dUa/kNE3x89SYBkU
C7owAJw744GrEdaNl4Vg8VN/FMdfHqAYFvM6I/BQPvIm1Pa+KJIW2p9fSmETclg5lQM8WR3Dnl7X
K9uTI9um7KE0yeErXVfWzDChfiTS4iFeK/RK+ssDt+ZfA1GU0TrTpe9NBI7mWD9CI/034vkT2+qM
u0WjYf4JLY2Nqg6EqS2bGRMFgw3HrOEOt8cWXvp5RfhfMy6gNYkaT4vpeohziLnQrHovIS13X+Yd
JHIiOyXUBUmfe7WcCoKOmKxWtzrX/LCGLHqu/znHW/Ui54DGpdbmnM5+arbhRQ+/X0nTljepdhov
zHUPERYdxoh1oiG+UIlYAQWPWKCvOlFFuXLn9z3clSE0X5LUkiavFexYGHf/8/bassAg0h3CnTh5
f3MRdVp8KJa/9QRWpVe9OQiKwT6rjPMPvAeSPKa3jPUH8V4XHHzdWN4nA6v++IEJfhXr7ZA3bRCD
rcB4hx0MeFEGUROK01iovZ3maHqk6RbJ17JQ85ioKytEF1BbjTgpAGelwRn25bF0dZ9qq9BZjorv
wYtdU7MA9tsDydhaUPdbOe7EW6OTmwTSQEEk0zAzmjzmMAi2kt1psoX82RC6/atGZSXs7rdKbDjX
dJuU93EDpey2ugqHSapJaHxPOexcl35waNoeECayNtUoym6dTuUhPbr4mu8lRU3wTS7t7UW3qO9w
GsJKwdpaH1FgldJIVF/zYAVXBjvCvlpjC64uqCEZOOT7jkL2RczcE/iVfIX1oxgOZKnC5uSRN21p
9PvGaTfIASac8dSq/6cSnNK+s2X+dcnCCDZ+wR2LN5evdHRJ32m2W1l91DFx7r8w1PFkJg/dBrfi
v6LiETnaHZ/+ocj20ImWauqbGf8cC/eCsAZRd/dewTYjVTYWV4JDlk0DKsWsxoBOTRX5n4MSZReB
ZYCIggGGN7hLgG78a8YoH28l9ngn95cZLVD2T1fPJnTSTlNhHYHgq86PbbYS3r+K7J2I/Lcx5Fe5
GW11xoFQV8W8jHPmjHDqv7dovQ5PvlKZP0BrAdOiJz4TCw2Lih45V2u0NXEC7ScdC+0PG4th+TAD
nuHas+bc+fLvf0HIpvezsePEvgZnSsap1vgCv/+RajklrlQS10daUh5wPZYv0t3ZSbFPSefiyfOl
H8SC/yNGMRoZSkxpJBbYPM5ATGwP4SNwJOEV/FDqoxfO3VRMI319JGKvPZ/3Aj9D3VUrVkAVdG/G
7tVwKI6VXkKm2bV2AXGkEj9p2J5BDuBHoID0QsgV9QAlWVKgMf+FzE+VeBia8HtxpR5+yV4OAtWk
uNaLRQzimQbzpAVk1/D1z1P7zaTU0uhJ+aCubCKUbj19QYQZSUlPQGOJ24J1fMnSlku653yKPWcf
VW75PAj6/RZCx0016zjM/Yyi1Ccz9oTiq2o+rPtQw7WExcWeWNlNW1SJc2JtwtZix/D2AhaGKET7
OPfexnMBI8a/iYDYA1cJpOKbx+gVyoVkuTO5kNDqxX6cTWi4oenSUpWlLldBwpqhrIshWYYZ3Zu+
7YdVTVUrm5GKMG6IXDY4a0Msn7AoOTqg8/ncIie3zbTXpiky1a28AP3En4raKi6Asc4dAoM693+u
PtlVzLdjfLToP87EsBPSMT2/AVJ4NfWe/rT0fFRZGK2W2smPrXYWjAEcMPv7TrU34IijkD+tg2cN
HfMvI2g1Clq5WqW+oOYJvTDLW8JFek5GvVzNXf5fLDU8DM/Y4a97sXr8neL+rxMxzSgfZNi66pRv
ropMncM83mG7HVeGV0XGLwqzRtPr7YipOKiULRO89cppDhYONlALVO0vl9tmuliLDSmsTSHX6VxH
G3xYL/w65v4MF0Nsc7iH5GWo83co6sVEQPpLUkvWcjk0ljbVQvsR7sHQAmiJvhnE/XWbDWHtaNb/
3K+fE3S1LRgK4jZEphiMRikT2rG2KFHrc5nhZTyqaf0dbq5ZQgdBggYvr+0PrtqnPUfdPqrnzvqd
W0vOdNFdOkP/altb0qYcFtl9DPiD9UQ0XKx59bd3zJbryzlnUbu/Fn7eexhFmqMqVYef1g4uovVd
tBB58PsVrSe5O6XQwAcc/mFA8ZE9w1LxY/fORM/URZDAydpqN8PRjwzv4fcvwKG/DUzmacwtdAgO
Hj0Rk9cEfXVeyvvgDJhajPcAi0lujPy3cOraXtGPyvxHcul8173xKAwWyfrAvSc5KnyUzOsBRFTt
Pwh5OpH1iBvnZGRyWg+Q9pCYk6ZVv1oOf4TvIXyn07AwTkiFk5Lmg+9XFDYnxcQrbUBzsWCthyHk
+zXO46NOA64F1PQapetX+9TYDUb2e0+o02qrGiVY/ATe87Q532AwezYLExzNJbSZu7rVoavnfFxc
i8IQ+5RH7x5XM4C11aD/C4ACdyN2FGsI28e3eQU6IjEKkcbChvjg2CuYyisA4PZlkAGHKnWGfU2/
Gdh3gny+3/yueNXSzYscy33I4S1iNrF5DGDF8dCkhePeeiojDTHfR2WSSmSZkRmeJuO3ZQtvosQU
1NDYwh5Pdcso58skJoaCuoEXnObqFOGa75DYdoiqC9XrMrgUyJe8RjZNUznDBmrQPh1xmTzYozoW
+cgoYXdF6zhFORw5NplTVs9ixQZI7/1jd+AvOu5EWrNbT2Gcf/4z0Psik2xHBQfVwqC7BACxPIV+
87+e8UD4hmJiKAyw9OTeHZIJG0hmOnPt5t6b/w2Ndjl/y/yjN5fCsTArPOIrUIuCpQ4S+x2wsNsk
+2WJNiFJ8haEIupMtamnXDxs/gnbLRbRWyhurWhO+iHhzgW5o7ElTBu+O6ZxyWTQI61uV5FRG29m
9S07g5RZls9GNuQSkKylgX8e6P2J0OnhCJkwAk2QsKUPL0UM48iiVLhIQUsNn/MLWw8zqaEMBWZS
53nfN0gcu+eN2xXKQEkhd2/lMWDW7mKkAR6AlFAUC1kSa7EDHdUhFZX89MWuE217z5pHRg2W7Xej
NmfsxymucfKydotkq/DXMfgcGsuP/hEiSpYdhsQ88ywFyQRqMpXBKHU8QH6/DbhmKtRiqu5z2Wga
MvGNnz1v4laV1RYpOgqSLEtU5F85cybpgTcXVk82xUoI9chP0puxqQCDLkkK0NvnOnwZI9XuyDuK
ww7/xVwLm+pKc/09CVvciwsreh+XiFJvk4o42UYa1a3WGl2AbhlF57BrUr49DqrVuvj3GSMm2xaT
ksTroB0AmBhgh31/L/fF0vRfEgHeY6d5SqQoi69LLTjRscEORRTM31Xky5vG/4s3ExWpAF8n0AA2
G4DcucrQhrpRkOH6Z+ROSxFInfvN34fXb6nsjPZ4u1n0LQtm9ML9o8T0m7XNXAfzKcrmKJRG5ZCS
Z9hzpJ4Px+OdugorAm0pULgMheyk2mRsDnHh5wKeKTaIIZHv/aLSI3PUXfpVLaHY9ESxrTFGrPhp
NAQVhxkwTmkVbb06e0JTW6f6k2QrkLH9SJOSZ2d0lUnJpsNA/IhpUkz8XfGDnfwk09NDeaCY7ZJQ
LqEyuiMJAnTvq0ocwSYug/rTCyMw0DPoyEbWdNkSSrd2N18XQdqxuTC6fTXlrX/Di0dvBPFiqldS
0fBXikO8iUpzssH6mxboosIVFCe/u7rlvmNJINSj3+YDfJJqX38+CiKMQjAJMiBrG5gz7/hWnyI2
bmdX/i8En3rjzW3wmhkJ8X6OtMSqW3rMnYZe4p/59b4cs/21vf7rg/qv2qMm7ueG2aRyD94NZb36
TWwJmJxE9oEaPlO18hk++6bq0JZSTLvnbQdbPmsK8JSaRpt4E231Ali/rsF7Mim8Byo3yK86Nm2z
tcOXafcDLOrBImwMBuZsHY0qKig/m0yFWMvI3hmsOhLy5TMue7dVxcqyB5kI3K6r39GLYDsnGDzx
CGgMSXBDDgZ5VcibEeH1af41XSxehPN0iF6MQxQ9jkie6+FmmVoHu1BDeMW+MYTn7aT8FjWr6N20
oy1PKnfF2+CPjS6zV7CGZqcg+btA3eLxGIVbI0wHg1vy1PmNLrNHSDKKVCRXVEvv6bMDk9rLioZQ
oFoLQOVyZWrtnWwnolheGzxwbfyZCaPdcY1oL3DezyrzsDDN0X1JuphkQA+uWYSZBHIKXIRoRAey
gSYN/4DhpUwWdIZQGOisCl2cTzIExKa5d8uy8CKPSYO7NTMw2IX4Z+TFB6LwxvkEFMkQuWb31Cay
wAz50de4//AXM0q/AZXBOteCI0cUVIJr5RrVes19Br1FcOHmpUjDZgDewETGf6JHj8lQ20Cjg5dw
4szbAOTb5mFVint3G3N/5lq4m+KmEnnQDInNCEfpRq2120k3uPG/qG95nngG5Z4tNpr+NUL55n/d
a9aKPd45kg9MsBT2z6t9ECwaPFMA8yBmaWVkOb2qS0TaUqLxEXUNpuHBw9tvoNCW/7jW6uGeszwv
3yR/UCBfhvdTYxYpufUJdGlp5kKMS5srA48Hrp5kg3BJLViLEANDuwsnoa/ci8Z158iVnhtLvekk
ewe8EPt5jxiSQkJ7WnxCsvfg8CAnRaTySLMfoJXK0srogqcVBSwBRwuQQnnPaCEo8T+6L59uuaLy
+ZODS1YnHNIU0GOlGa3QeVnR9gslxjVTE4qYyJjz2wAoFn6hKBYJHOpZf9+tn8KOPv0yht81My+b
G7CA+Nrn3W+EL5sh4K9neagC2t8sOHo79CglWRD3X1wzfaY+0zlhDPS/sshqj3s5JF9Yt3YqkmBV
5PHVyGwXvVHyuptWow4m1MWUbpzod5FR0kl/pQW4XdoQXoO69rpc6FSwNm2WnW512lGEjdGK1ZNu
dplpPNcpDaWB7Q4HWat8dp5XuPUgaEmkrAOKzrf0YMRrcSCKbZ1eKme1y5hwPgP2Qrn6KhUAFOkV
n70urPclQvSJGhgEcC3Ap5ilr2jGDQMYxpEgcEMldHp0Ndei105pUblaxEwfJn4/HWbUi46ikSti
K8cBYqL9ANUrfsd3fyg6g18qoNENitwqwUdqeOXmUwJuJ8hdb2D8Lg4dGleytib1NT/0p3AL6yT4
ZPT837awOh05itHzRI7FM1d7K0Ti8qxkJI5Mx4YhjFKq58PKebK+WErpS/5q92XLeHZxq9Gtkr4T
E9HIAwfO8B0LWhhJ/bz6V7KyfNAr7z/1Skmrgcox0f8FrHHFRECg+ECBLqJSpmodoXiwQBn28Aij
+O2abhTxgGrqaRi7FkbmbNkF0Y0i+07y2X1yiBzHVA7Vqol8d67oLP8/YZQNHNjpt16FWUcN75cj
5M4u41MndweL5C1ZA1yKU8gnQIY2sCPCQ5IesbvL7etN/G/7g29FPsY3oJx3Kd0hvJZhEcsOmuLz
289kMIaalCRJht+wvADfMlnKTdIEunq0q3r/QcQzrR2M+FP1S+c60WkFAmMZNiVxAMpoNj/dZE/C
VSLlku+QtH6Krgue11NXgPlamfqV3gbHycRyK4BagUefsuKYVdlSJ9JVY1UAm2F6rbmnwcE+JYyf
DcUFOcoMlFE8Tj/1DQBz16Uxa6Fwoa2n0+Tz4vN2XPhQXwS+VoBAiZUMM3t+lmjVQBoagpHqYUM1
FE5M94meFQzqC1rwipvRDoLd+wEbnsjY10+xZR7cxhYg3yddumIKaW8TS++ykxqFft4/t2YGtPmN
uNvzDtzYVKrXGvKLpuX8MEcHA9hVeyNJdGPN8mMyCg5oBgOjSZ5xW1y2b5XF4OSy4vROhZWAjwB2
v2M1JM/KY2EhJFSaRiNokNVVcdpMkl1S0MfmicWesLIKdpU+nhXl7Xf37zLeEV5yn6rupP8zMs3L
e+DYIB6pnuDR7nhslTqbWzmEDWS2guFOu/4bnDtiEuRro3Je4FsDKib8vB2P0uhST2JK2pzu3HQr
pJF85bCs8XhTA1hFG15yAfveWaBZslDz/YqAFOcFKUTjU7gIQKrnG/ROsAZcmBtKcxBOQPEC3xXv
Gu8bN3SCqH4z7zNn7wJpMRFQGHSlghiy7CyfEppHO+p+1YWtW6YnIN9QKq4jVlRIj1EIGCDotZbd
W8H/9URA7tDVEJXjSbcY9b5OTKASHSl/xdaT8GySl+sU8ej2A9ok1ml8maStScW4Fd8fUDwxot4m
9VscHc2Onl9J3HUXjuY8gZz2iAhs2tlv81i7PXfycKPYxvr8qjwyGNfGeQnWJVqfyvSbeZ3FoPcw
2vnCtHMsZxMTCu0a6jLUGSjpwGR3bBzI6QTI6iwa2oxf9N90amSn5Gm3UrQk6YWyykN1muu3IFrQ
6cPEKcaxBmkcwRVLwSmSdYlXCc9MKfGlvkBknvIpxJsp3rwtfvK/RUVSYULJ1eItXpJmtUfQNw2y
lEvYCWUOKfJOl8T4HwblZe58YzsYZvbVmuh1AzZV07GbmxxxtRQyjt24uAjHm+IH02zeju/UTK7s
xXIN5psxuuOOihIDMpmZW2Lz56RhZPFZ+8a8xBiTZMYetZnQhh9K7OwCl04StmDvwCOSWyfULQIQ
9B0auQFesTtCoLnOKs/NKlCzG/z8szQDRiccw/w7qwqOYeGyg8hyD3++ebj8h0Zs9Up0TeItZ4E2
JQ1nw0EZGcb2UWVubO9Ti9t/pu48ZdDLxqKRV3swcwWWzi9zPQUQzjgbzk9rL6cLKB09/BKz9hwW
4KnVpt83hyKqlPw7lQMMg/BGJ2PrH/X/9hXuo33yq5fmYB2Uexmvuh438LB7OJP2kPnbAmWcxIkv
R74vFaFgcfl2j+z2W5i/ZYUZ0JhG2u5uVhvFmOORvvqYeaFSZtqRTjyufDj+EtmZQGlfAttiQORB
NhhHAI4Zz6CiztElfjwxMmn/4nO90T8JubDRaFBN4dA308QkJSpBQFm+C730p8tEZ1/hkREmZc9G
DA+I7aEh8+mVOhMDlTISZXiQDcvZxVrJURlTJaAfLoiruD493iQDkiixYRRqBEmYGXOI7PZtmaGa
yEiOiTjvS1mzoEjOR8AlBDi/OvDWFgwPyWWl6wKuyKDfdkZc8mKeyU64/FAnaqlrHf2c5Ydl4iaM
qTR8XInJKZTHkUSNP/anHmg8dtysCmVmio1d5qAYYUPhwuFycG9NAGHinORLLjMGp/puKydEoug0
mWrkOwKVuYORoZNiyWIp4d5ZwFr2ezqzuhcjLHtnaYeorImmBE2zfLhxkpPGMJX7OMm5bep4dKNo
o+QHXbeXnv4K/K9QkYOzNkl9j4Ed0Yu9/dSB686a1FWcX6DsMx7fXFMu1TwMGHy/eCQD7NqiWEzP
FHkB/BzICLbdnnNOIFbN4QxQebI/h2ktxoInqMSpz7JCYGtHuzlDsI3cPpAF6FC9DzKAvkTKZ5Hs
NmD8JB2wxnkggVcd8iwTXya8C1CtMQjnORfA99WTGJJqRN3WirvCiMNSmpUVLDHVWHqjOWO6FRlW
WpQeZhQYLdvjA8eKyMY27zujgQKjcVfVRRInf7j1ibBSEzo2gYS9Rl++oayvex/AMyFMHPPpBvHe
g0Y8fj+da3NrRpG6AF4WKpvEoQs8jf4w+QvBw5UD5xQZCqXrGW5zgVbjKJuovvqRSiTIiUp2AIec
jbeUTJAKK2FgcyQEbhaEEs9I+FEUm1ziCHBkjnrJ/2VVSYlTOqPr8hOLf3mVmPQp9WJfiYdEP9G1
TVpWQvJwT4XylgL4eyz93Osqd+WdR2qpU2wNtPrH2SwFfFYWw7coRgyWSwTCHx4/ND+B7z663IUG
xpaOYTh/6F3ju4VrZs7salFSyxSZJNxAxwGqScQpG4UfMK+4HbT6vDyvK4kJaZLM67ttQN66C9Lk
/Boj7mlpNP/excDMSA7tzIuRyUm+FhNcpautFcFSDnlcUgMh693FqXZtCAuisEptYDv6M40ER7y1
JA0X8n3qiT5+Ik7jbGkwvBP2E3kNrPqqq4V1C92KgHFjXYwiVa0w2JMv1O72XFlZZqlZL0/hPHIN
1FLM8PG6k+fKsVrVjYq9V4KDqR2ve9IEgdC8S4z0rFBXpBkbDM1bkD6LSYU5ljjAewth85vSqrD+
SS2hdr1tnU7VynejjwDJQihJXHMv012aTid8ATmjs1RZjmN2B31SpWgA2Rh2EzbNdkJymzJBvw/c
xbya1qN4XA+AIO/JDFU0/edD7GPtZTPU1BqtK67Xvt7UdeI4sZMfMD/RS+6lpFvJOLZmApCuroK5
8xg4bDXyNnlav2ZrjUTobx7WnPFGQhV7JwYVztVf7/Le4XJ/eolgkgyYfZtWAI6tm9WnK0ceHC7l
FYk7SQCQRJvAWGerjl5fU8oX9tcnPPtVntamwjnLxNJF4obneaCA82TXNdRqVVgb9y3yLmqEBS7L
bp0ep7K1imDMixBwBd7qJy0HzMCjrN2HHdOk7/StUZfw266fEw7ShNmamVnMJclzFHDTQsB4AJJU
zV0cM/0hSEZxuSU6Ns3bSt/fBMNzkoc27V0hWAlS+Vexs98obSqtG3gChTA4tPFfqgc36GeaRDgN
38BqzEV/yuZpeAO4WA9bufB5gyVet+9dS/BG+NbfUWTE9onKdKvBCw2SEtSbN749CUSkXIMuU1M7
C2uHJPkYkXuYb/Jq81eOKf3dax2zicQCjRhDdBAwoLOR8kL8kVaHXwBP6GzPHZQ1yFFc4JQABoaJ
IDGv6F+kDMmnDNbN91kHrd3Q3NEmZ87wvFFWrTKjrPs+WQxyM5zu5nYZ0Fu/R2jI+wMwPSAqPQid
aRDC3wTc4gloyRsGVH/CtqMIYZCJ6lEXnFPh25nHPJs0MhkdGZ/husJ5s6dv3SE+dKdf6H+CPd23
Tar4/P8F1FT2NoRK8jzRCYu2rxZ/lDZ8kmm8DXUBgX0aKishXg1vTH6CFvvmDeGsHUhsurJvrqT0
87Eu6Qr+0v0ls0lAECSkuh7veUUiEo+6bPByCIRb95LsvW/7jCAuB8nj32rcJkzyO9yeYxo9tZJA
kjT8YjaX9x2lTFLNjO9WKbCjLKghC1GsOosBFAvYUSVHVn93UQxi+7CM8ZkIdrKRGVSGWOmdEyyD
I++M9y6lwR2EoCGLMUNcQNw06E2B0NW2wn1BnVNFK09nOGFs4M4VVlOJD0YctdeXmD30cIosF61d
jN294m7iiR8Gh3jx+vW8rxKRMJ6euWn7hFDicKMY6qZb1xFzqBdfdwNhP+KvIJ9CTGPTq5YebMqN
dbKU7NQQuv9FQKuWcXwke5QoXlaNiqKh4jscCJfezLulPuewGfZ67g3a0zuCFgFcuCzpgs3IIZ+v
EB2XgGDgJVeOqiuEx/AKBgZ7TWufG+rzeKhppXYKNBLQnGAyhtswIz6LSCDTC4V9FrfWmDZa3Bsx
cbyEeuLKG4UNi7aE94IzxQfWisQ6PTrdSIQXyvFN8GROTp0NjBV2uHQeDc2+/nOFmlRtJWACBFHi
zxn43cr7tqIvbMLVqmgbeKV4FHmm8acUAqre6DPvNYEbSdg1prR8bw9EzgjgbiX3Dbj3n1xuKpnZ
OWN/vorNqSq1IEIX+GXaWWddU4f1DOj1MiBoueiAjmDOz4ubuO6/J6koUz/7jHhsVU2hbOyhopWj
gc5B0E2fIkCFhr8HfKTYwGA6pOZwoMkGUgmkUb3TH0HoIG8dH/ezVLG9/o7gLjv1v/JSe78jBpsz
DJwQrHHBVIK4ZLK++e/3w2TWHAzrw8grb+0KyjeNZ/CtQvKs8E49QpIUXOF31F3SVMD6XATJy7b+
P9SsyblgMH2rFoCnvuqNKTGNKRll2N8xdgYl3tE0JxT+siCHYFSC+THJzcS3ZUw+syp/Koyc6nlf
FA2sKVmW/3nlTTk6D3cWy8p+p8OswkM7nuyLf6rZlPlpt5D1cEuJzeOiyG0XQI9dT2hVlKuT/waz
Mw26E8by+R1FQgyVj0JE9CPiRaI2SYycNzd81kasHY/DjxGsldRTeTjtPicFl8xO8RQzvxnDW/e7
zwq3xogL3n8fLAdjSYDqvNVfperqNwPdmQ2qi80Xn8/13oCUqR9b9SqZtEO8UGtJtK8ALHESRbzA
cJ67jv8cw0QENB/2N4KLrG8V9acOP7l728AojXFrLZa/j8cSnnutxEpjhS/xBgroM4a7xcZAiWPx
tHfA4zjxDLQFMV/kq0VVRZcfOqcNybyi156qnwcZkVWbphAyhG2OeePU42za9yX7Y2iGFhMdDKY1
lAVM6QEKERZMRGb52Zp+x5risdL68mWW5riQTpCPO0UAEIjvgYrhxDH9DlIPb9oFDeVJcYDKg/K3
qBhPEQTUyvPKxc5SKct02LQxu/1qbUVkwwHbYNJxGYMMBlZINOTRAByCBihn45398yNKwEJvnQbn
OB9l+Sz0lRKth/HTbBqJcEyEwmnMmZR74bROVG9sL5vQmfxN172xtUUjNLTqXv5oKD4f9Ty5oQLp
KRtnue0RN44W3eZ1Qjomtpxzn89AZhCwOq/s3qBlk1ITGz20f0VeGeVmUFN/auwEldiC56QrqiSe
uH5Irkncq+AtCFxBvxkv4AUdBoVLBIV5JIBCmCpzlGMD/b4o53UuaUylhMbW9JXY/OMFykyrcbQN
+zhJ2sb11+RhRHdzUqy78cpTFbTFhPEJD/B2+yBBZXYnNziPpDG/cG4MdOf+kgSNrqLulgZafvDq
eR1hv3cMgbpepofnTsKKY1JmgF3dnxyMrIOwls+Lxdxs319t/tKS362kKGkCivtfay1hLo/5uZss
VTnCEIVNmO9TJOtehKy5guSnCX+nYQbML3DqpYTZY9yVBW0NDCk/2ZThoQn0GkfgmY4trpkswNQ4
ftrG36iaHujhft0sxR2OkjVfMw0lJsSWd/N9IuMoykBx4U/sWmtZfv0Jwjt+fddideein41bbd+a
GyOzvDU5P9Ob2JFVuMJOD2vGg3oaXdg0HK5J2suphVN59fOMRMQFZPDCvkKBff2gnONkC//ZPU0u
sUSrh7QDssg/Ek1+uAbZLMBHDMFPjSyTA6JwNtfn3nNX6Kc1H34UURqgfVq9/Q1wX8PP2zPUHl20
566vS3rOrpi3AgNSGcgmQYBa+YBKO3TS5H8Ide4VF/JTH9da0DkzbDB4msJyvZtfu/m4BBqxZmaM
fLakWUgZxlwa/xSundDY9KsYBecLnot3enq8KKXuHin/SeXlYo0gVEsV5+t1qyMDQ4My+hJeoqvr
1hZCkuc9AQqx0jDozzmao3GiYl+NZfUKlSGnv729faHwATonjb37UxinQnTMMzHI7wODtUS+2dYe
Ynzd16sfcXxmnGZ+AkP+fqgTidwZTm1X7RnMAueX3qOedDXJIW0hFU7DWCAF6mlQhunJh7pUieQ3
tMvGXR89yI96/vVHGbCcLdArFSAY0RkjktoiM4XC6QnR+sjgTlgL3fVH9HBVhFVZtPLrIS/QPfEO
GLGcOOjIL8VZIfdZPA6zS1OP3lJsAKd4MT6+ddcaRO+VnG8/R6xGPDnqVyEbklq5TXiZw6EDShn4
iI9NqmpZ+/Fx2QbE6Zgi1FxYhh2xPnDrQ5XQU1zTnlwyi1BAbVhRZOThtpmhCZWGBgITLEEi2kHc
g5/BYx2RQLb1myB2SA8pRuM/O2wG6JugFDZf4GM/egs7HoXgEGBae7dr+YSE9+ynOp+BKcom25FH
Mg+AY5ROeAQ2/KdKMeUcxl2nYZ+MdqfKDgLXMcqU6ZpHu/IQGbISW+VTnhsJvwncGzJh7Lov5hqR
YEKaMHy/z9En5Dr0tI+Vm1R75KfvQrL5zFhkllrg/zeJbHV4R+uN0B9SkwbqfYUrhdXySqZ5PMo6
e2NqiWdPD1eUCAUcX+E9CeI3SwuAHcNyn/LFhyGODrAS73EFkHFPztDQvVmgM4iKo3hzcvzH3i2g
jsaWcsHS14H3dF7qLUqe5TK2O6T6lk6fmX/2H3K44RxB+xV694mBWetNVxf1o+yXN3O23gPHILUp
byAm+J6rC5MRk4GZRjz2yKz7twBH/WDQx2ghqOpb0WRDfAQZMZWEcmHUsByjpjfya7inphx/0Uw7
xglhxrcD/JzIZ8MNzAORQdrpfBGxzDok9DfKR5JLbsjmmnAkPk7yUMPfR4Fz7+U35azijnbk7I1B
H0hRIakUqM3HRShMrTF34LdZypIa24ImtxlRzuSTOq4O7fr6+gcyl+a0BtYFV3anL6FdE7UChFGu
wDl2o3X6s3bRfedIgHQBBG8EZWlEiMbQFg8nsNBgKkCi6Hdtspf9LBwet33JKouqx1wNHCnym5Ly
M1Q0MDdcdGBFhi39WhtWtoFPfsWeKwZhvQnnMMpSTkoBiHvZWTmxSsXUWEpKPp1F3m6DD8vwcowy
Akt8LkQbYUFGdz7Vu1YveohQUKztoZu52hJtOYWHO108XsqcfmHNKt0BuQcVmhBmHuiaWfR82K1V
SCpCZ7ClkYn9S0HA+OajxF4ur/7PYxppFnTI7GKcnbbf8+B/SIaF7fD09faVsUTosJ/Va640VHGP
YedG3HQgXOU+YGI32l7BzlHWnIne3CcyW9nfDgpZgQm9KvXCc9eIKRjZPzjfJEhQcGlSss5aap5t
gvn3QLN/9kyGOjWlPH2zjlXd/unqDzH6JDpU6S1RSHKQUP9+Zv2vY5UBA8taLAG9iUYiYZmd3iwQ
xdxGxCX1QxKbShwq/8V1JHMfkujOPRsVCjYALAv93iE68bWbtDStp7y3aHADEQcx/g2Qgkax2k8E
yzWOcDmbUDDkleEBPlEe363cnEP3Ru92F0vqw8pzbQcQoKew8DldxAl9Bhl4fF5n+lJAiddVnIVv
fHGV/Rv6vOsdZKi9FweTUlwi/r4UQZAVshhHR6iHd3yMTPtqZSdrZ34ulSpoU1tYGC8XxaRs3tBP
1ga+hyvIWpJlQUuGTdY38/ri4oUgnLXj2TF0PeWUC31vIEYLheZ7BziyPgaa3112po1WXQyi0sMd
bLmLHh11UjmUtWaboX20rG8tffiyyiWdA89zUsnRmMLy7rGAWCUW/p5HNZ6IQQ459FbRPWSa1KKo
kaS92AvkojtKbSZqjx4W8yrH4s6wxTaAdAXIZS4Z3VaKIpBJK2dDjNB5j2n5jwqsIxmA1t60kVUL
28fOk3oU/QYuvvkcX91ggXcipp5efIivsJIb1Utqn3RtVUmUM3R7MmPT6VevcilK/n1KvxH2YzmB
D1zgeVeJ+zXodampB2qUGz+U6VYPPeS9j+iy+VicpkSdwjoawHhgyKcMQRYMJP54Wl/hcmOsqf4F
/j3gICFqlCnx+4k811jYOYyCKRDNTqnj11FvgFJO7qDz2bKbyOnQW1SKNxcmB1TFHopUx5YdZjop
Yh36Ltv3hsqpr2sBux8uXxXLbfYkXpnNLLPwIqbvZs+ZHpNb2urqZRXKV9ZxoSZeF6rHMDSW0qF2
583XIAG66fYu5vbwD4t9j9APPkq2HbW3DDo7YKqEcZ2CEdPxsd6n04A8cZaRaWKOq9dtyKzL7iu5
Us7oWmqLWMJgPHTngYIKhcbP68OAWpaiuaP5K3VvG0Z3w+p8hUeIQ5vJWXMq5GXbRw+O4H/HIeEG
jEAbr012ELyWRGDMQtYdfc04NCUwh375c1j8J+jpRr7QtIC9EuuoJj5p7jFfTbEkoLk25Z5DZ7/Y
S5PEOz0Z7hoSJpeoFzP+Gjn06Ks3bHjIPi/TKn6AwsAZHwWuDVpa6pLhmx4tU7uk+zEXkzDFvAo+
nxpe+LGnd6x5xbiiEOwOjaTD+iu3Imv1DTCRcyN+qhBasZBTXwO8OaJJeJE9IcoAHA4upHWBPPda
0rwEisvpPIwUKlm6ZSHFuNwnGBuxf+cNsFbk6syyxKhKj+7lw7vP3Drxy4SR6dmbBrPXxBhX7mED
7/7V3B9jqjlIhU7CvMRIRMcJ6unLfHDrrKdLiXHTKTHVzeR76vn92PgYYmoiyDCZ2qt+BmyGSez2
0f3dNVzoqYXBEU7L3W9QOON9tEm2eccWGQ7KgMGMxfp5vNKfL9dni43Fo0w5kMd99A4R+IsgQVj1
kfpnoXVSiyMUvbxUhB+KaSSOBOSO3gwzrU3vf3Qb1E9NYGQjqjfKA6FsX2LugT/9gA5n/O3HDCGh
ehkZInZFO9afr+axmoXZax0qA8bLm0HtlrWblPVaQNRfJzQ+yqFnnaNrYCQqM130ibWYfLKHpXvn
Oixl5eQVcVU0zm5NCF7kdTeYJ70vny2cTDVV29jkZjIbCHLCz7U8jf9zySydrn8cmYEA0/OAFUe1
CeYF4GuMI9JUl5YrU5b47UN+7flDpeZpbczrsSNVy+NB7+ZVWNnwOqyC89hT0fht4h7UzliLivii
AXlIgac65sqBHtB/PvgxdR8yB6Vk3ObYaBfPZ19AgJLJX2KpvGGdfiIYOHWrCOitNUDLU8dlZYYQ
D2jG0ZpIz/OB+FyvXZ5Gm9wGtt5mm1RvMdMLqhveMmQ/ms3WjAt70j68gUF4C8qv/6xjrIlZ77w1
P713Imn2uWWwWumKS9qk+rOLaXmIUXOD9davnNtIgg30WgqZP3pIcYDsqGc3omo2Bn9PV3CHyTU/
43gR9q1S8LKeQKFDz+onCEiDeyRXos24kz0/+o9wxRilC2shGm7InjmUaY35CnQ57PH7kjNa/1pc
9XwR/nFIJQwyg/rAh7plqmmVjAEXYPWxSarQOXKnTFBSGyjopEHPKwEJvmmHuhQBKDBAVazyh36v
Bv3Qpium7qUhIpwOaj1R13oCJN9nGkCPir705DT/k1isQrG9shJQUsiE6+I2S7eGbGfYJAK33Bdu
n3R7O/6+ZyUt3Z+l+D0VWWCaIfANZh7CHnQcM+cymMpr6F+S7jxgNRcECI9LraNGULqw0oELn23u
D/mV4CLv+VgmTQwGJGSfc0LG291U6Cw3iABtf8EmZRwwqvG03pcsJ2rYY9Bbdpzi7/RsUx8VD1As
mxqf4O735xq6PjKCOvn7+ePqyhds+JR9uBsQBUTqnL310kYkefkZY7fMupqP9XhPkTHyIKjC4E6U
SUW0AjXvGxTRDtkQjrlADJO6amLO+Cen4qnTQS6+h32tDAJSdq/hNiJ6puoFMFHztJUeBOXsz1uV
TXhBeSh6rvMth0KE/Iw4N0MXKv3L+gUYkbz0+ApKLWuXr4XkrMSGgNo/ZnynmXz0Dh4lgY7lLhV3
OkF/kAg7o6nGWTVQ4i0er/UrqCxbMkBtROIc03R34Jm0SVuWFPeX34FfAVw6VJB5KtWVcPVpBBME
ySxXY17ifJMEyiDB7XLBurCGT/bSRmvW0p2fKX+pnDF6CHsxx7YAx4XMde9VsLXMvXQBki31HWFR
53kJpV5unyjWJ8rHTBqNPLt7fIzjoRmNocXoPR9B76aBVepcIJSBIu3WHQjTUmMqWw3Ket8yjb+1
Rv+sr8qmnyYpgEMDUCqqJyV9Wict9DbADXKwY9PqZY7BkFAlloEgxKwdIEa4MVppcAScjndZseMi
1p7lPyJwtMucvTEB4viDGfFSj7AgOIKAlQL2msU2QWWdx0CjT1RsmMVYNQDaSPXMOdsxobHhly31
UuwGZoqLX+6som2wH5WXCENwXmaF9EB8pqZJQJXXvhrP2Pu5PVzNc+5RocNtW4LZ22zHbhPmJY7h
aXJu0nL4hSgIiUwe4z4wlRjmp3zLw3pELgQ60RQ5FU9wAFW162tLdEmvL6Kpaan7l6eXLOHqg60i
s/ql/Ni9fGxIgNfg1lNpHFI0uLUMTUCln6U1Ol9ZlHI9iPdJ6NEAwaAuTIgVTuZ88vRPxkr7Mncz
gV0hKKy6CnaprCaTWl0ZdFOaEoIDsdYi77/3tQ68hHyDZGwu/I5lt4XkB+D0WuE1nxRki0Y7Alai
46+mNrKdJaG4dcbWJqSkzwUZq2loNAZcH1Dw0uhm51wF6MsCA/mSwAXiphNUG67OBChiwRiRb06y
7XPbwY7CYugxPGB1adaQEvWTqvM660wayGiEPoXdvt5E4I3N/pDcpTvM3v8vF6+nulL+SlaLF//f
d9kakonUH41ob1EAPm6A9T9rn9Smrc/YNZuWIgCJOQeDrKKW4DN1J3fqLMvbp6XeOpQMdPp4F+WH
U9pMl6qQKZLivAiNAlFyTSu4Dj31ef05il3QomrY8DD1FjWXa4JwhdhB0ZJSTYrN0kPytfmL7iVI
j2FVl8GTvdvLS3tT3jMMUbSP2kNgFthQxGWbJ+4MoH7CiMz4dePCLUpx2NkzPyTzaiWsf9ckrTaN
sRP8RQyvVkBBlkNaE7hgyN53luB54ppxgkBt+zqCxbG3srInuJ/TTNDi4FQZu0VYMB/jAbG1UghD
da5XpgyRS9UJZCu0/jiNToDVWaiIjEyNPr3PcuoqI0m0CMkSYe/GyOyirHWwK5BAC5h/RBgntEq0
GGVx68oYrd29zjzD+Ax40yseiZi06oA1Y4r4EOI9dQ7zBJR7OBUHk7PnsRwUeqx4yGLZ7kFFed92
wsRMnmMR05EaSWzjdA6CaSYwuAPax0SqG8zKYs6rTOZNMROCbH3i7SGXcBRXfCeCTSh5y5Ku1zH7
h3dtLlFrglTuZqhHpJfxHJkYNSMbATACC9N/LvgFj7de6GqIAR4e+sto+2kP/Jxqm4byNzKAmBm9
9nojYTc/nC2paZR19+cidjgjwjNL8IX7D47aU+plhms5Chis8dnQC6bMIWNg3FLhr1h+2n70Z/zh
HgGwpQc49DZm+XQU7Q38M5sN5ezC1Z22mtmFHAG0Sz+pp7skG6zXXrPJGTPQb98VmMGXTwZBmBK6
53ZF1WcXIjxMmMbqFYO3/MJsf1CDdnhBXhYusLNgfy+xPUNrXucRHDh6MA4CpkND55hlpP/YVlCl
f5InolarzvDAKuVNHH6ku2kzkKseidwO/nrX3w51ymfTYdU9Z7n3N9DwNWECXRIFLXd7TIsPU5ei
NgrBiz+NSmfZkOs4DvFCKlsnvV7RIW+07AnV63AHFXJkXByy8a1bl5zCcqKAJTTjRG4IiR2WQPWz
uYnE3KFyOiVg7Kyjoh4svPDhzIu1xH48APr8xb1rB6ZbYALJtfEHBukicgBfnNEtI9bq4AqQZIwo
S1OAvCQPKIBx/qeC2N9WJEaiyHrndmgRVXZUvdk+Gx/F2pgOKjR6FaVOLaCOVtV2Rr4jAfTR/ryJ
VgnYLs0FPZzbak9l5B9K7eVcIyB1FMuNo1ABTrmvByBywXlXXJosBNN0WKqLBgtw6V8GYNt7dPCP
6CczQY6xy51fui0lVLghH0qAheJ9r5hkEJNOaCNIFmPZ1g6hunjgxI2an9NngpqsgBA9QLgNs3BZ
b8RF7R1IzQoIH31PV8ngjTgwP1GOuBh0dDj6oYDN/U8Mex3DAGN1qYn3JUl6I9kybLgU05G9LZUI
Yv6Ft4CQlDiUUfzBZg/b6TzV83lYOc4/caqk3hH7xQstOISb3OSaolyvMwHTy4tRM9f5bMSu5lMJ
TPEbsi7X/dPmiNgTrmzA6JgRHY/HlO27e26OySXQVcANRwF0Mgbsc+WGVCN5l8kYK9bFp1EnZZFb
8ZFPIjoukMWS38SNmIJUV+oHXTJ2pK7X9O5pf8FWM87RlCXbsBQ6uzz4lFUTRJiUG0KWKoHJBlb2
LtrtI17p/kKY83qnj9ajvmuTcRWozmKZxq2Xq1plkmwewyqw9TC9EUViX47OCMeXLrCYFUjMaI7L
LYjxTi6/Y0jgT2RfbH48Rv2zBhSElZEJ29LTeY2sUHMkk+hHg0NpH0D2G3XGgaUOHAL1+CGTUEz/
G51p+3thPkrm/6kIF3qJivQu1NIZf4aiQpv38Bf0bTmcPsKNd+NrKoRe8XOe7yd6O2ONeQfqdxsd
NLMaDvbzYjvPG/LHNwROzk7WpP05jeugmJKc0vjaQcTVdbfOppTxrvLtj2AArSES0GHQ1dT6mj0W
coPC/MoQ29iQ36rU8HdHizQ3eFlzQiK/ARVAQuJ+5zynzVFf8bg8Vx0RTs5ZW94rX5JuISOPeaTA
meG9QRH+4oZRnwWZ/g1hrA5EBjjE5Oco1H08E7/SyD5QOJNLyi/yaJ1ymvi6DbEqhJldIXQjxt1W
qJJvdhIwSx8isr/z/CGe5K4uFZIecQI0lAZXtU8uyUESUs47Q2o8+OS0kY+++cvQU2qisV2S78Rb
aQUFeacwdvl9zthsO9Fz5FdpTc070ry2lhLHf2c+beSe7rbOCYHyaat7F8LjF59OOD1LxOC4fsc7
dazpvaLH4+tBJTO1LJJXAeGjw28jzzztiUscC/c2L4Ii8KE0zwyqebhsBSDXMQxYqc1Kb1oLIzT9
WjMrlG73vFN70r90RbMzzt/FXZ0fKKQxQ+VjQD4PMnMJfwRevHpwFDSD9C54FmOtEktqsM7/F2tg
fCb96o0jF/ittkwKfHI0UC4J0fIl3Qr/lOsaU1481jc/aF66eBWb1AZ2uxDSn4VNP1pRgXL2sLak
shdkIevUivkSAATX6GSdCUT74wBSWQovtppKRSYv1nHUtYjXCCiel7SD1kzG7pkO7UD9QmTswWvO
JFP5T51Bky0/oJjp9euAu/15sCbmSDHkRUaLDq5QpbXcjn0tcT7UOYu227aBn7kWPXnCMUgkQqrt
rmJnnUf7LIjOBZGNUl0fz+dmeBOXR+MrvIHy7OWngvjham1Lfpixh0KDyJThkHL2JS3PHkUPPA9r
GVAqwMRFN+dG07HtlDBZafbTS4qfjqiOW/p2ggqi1HKp+UH0pwy0+Jti4xFE78SJmOxP9VEoJqnh
toPPfYw/5h8W/QacF+xnYSZU/AX+Q3rMHBy2NiLzim/XnKKrg+8zi1wjwBxH6/b6h/Af8u02RATK
ajjpM8lslkDeYqu/Wqu+K56RJ8KAuPyYLm3HS+WBiveOtWvmQSMNEX2QnKrZmhyQBTxN6cgpiJVb
tf9oda80L6KHTiKFMjYe0wtbVRrX2PEZPzkH9Y+A3s9Z+E3hkLJNZNwxjW2LBs0Mnk3Psaa7GGEy
w/p/g/LLScnvgavbAj7+ViYDBo3wx87ywyG/+QrVioREUlxNnsQkexQsAnZcLUiMBlHDgS1X7ILq
/Eop8MEt+MgRyOqfFylQ64UJjEJBc52oYUpAQl+57XUO/yBgqK5nv6HHxCPzOiiUQEQLdtdPg/K8
v4N4RS7ANR7aDFKehb9vqdDlcjV2zqNu5gwQaZdhOXZbnQB6Y0XyTHbNmiIcJemrlkY81i46pjAe
M47E7Rh0/sJNsflKL8Ns3nUfUTCIy2U+AEph7XY7hHMB5SOqI7cRI3mMxekfWUMMbJ9LEcP5FXFn
Mp5XtFeW7sAsk2kniKEvUSbqt5S8/T6YpdYc07xf/is8M0lpaoDBjxBuRcZ28nSZAwl/xjLUWbmQ
cyQZB2iHcdXNDYwqkOpxZoisp28K4pjCx9jiymn77rqS5zI0uFaRRej3TYyWknIbNY+oQDdg7bGL
X2PtXBcTZlBM/HZ308VPPjs8p1sGUoBlkaVzP/7rf63+7JGlsXnwkxaHMfVaWh2OVP3Vbmwq+YrW
Z9xPI6bXBF1/kRppQvvX30FCD51AS1X8n8RTu2IJOyIE8/qrh+iFmpmM/qmgbhBxqj+o26rkhUwk
1gSLWmOaiL4lqDhCUlF3nf+sV2cKFerf0O07ckBsyl31SkQEJYU9ufyVndfS+TO0dU3xKJ3/mmhD
3W/4cf0UkE/GMyP4sGVmh7sMt4I2ZFnNnlRu2hEbgZGLvx8aNOBQSc9p+6OB7+rWLMKWnUbRbSty
GloZcAmPmWy7yzw9KHAIgaLM3aS+MGY+VXqIc00LLFjI1EJHOPHS1sjyNzr+IPdbLCdQk97eUI3E
+WK6bxC71ichoNWo2exPFZyACtSbrO2YzfjH+wjx7cUGJ4+LowpXLG3jQJh97oynTU/GCneTYyS0
qO30pBfL4QVynr82wWAVSixMpiVbN8CaVPeFEnEByCZhRe3c/wdoc2I/siyKumsz5ChmuwFKlB4F
+eZ9fqygkQE2brIm1QlQDOFY8evrjmlk3NONU5ZUvf0t18ZX+Q5NrtPIBapGZG3hnKGxJH0rOYEj
jAro+wRiw0iI6jF2OeCwqumTa+Hn2FvqlGwtC+s+SqlfbeqYqJyQMEOf4YfPEErhVCFZMZYMOqBr
mmvXB9SlsHybsabzo7iSh4WoSaJBLdulxzJ0uTxUKN3COzSvM7NaJDqZL5OVFbiaa1oM5DX3xvP5
1aYAxlMSD+zPgGAv47qS9U+yR42/VBwoGS3gnYlD8UoCD1TNyXW6KaXng1kptQB9PLw+awI27bMG
toJu93AEMxzh8DROFiyH1X6S3DkQUlGkZc7WlTTRREuLyuovBwDijd5Ws/wv/lY/mirGwBwK5KjI
D2pRKaIr/PxLUDXdZe1dGR0yC5Tne1G2MdN3ONUJtQEo8QrwbwobWvyMG9tVZDpboZz3QW3BdKFy
weXxoKXoTCqZegzEuQ3vynUyFAn6ActIEMz3+jwADu4ot+idwvWnvwY61syWn2MhWHRd55QUAXud
RVLzg5n7JdA8Bj4gI3f1Tj9OTEqkFGmhBxu2y+ydfly4PUT6Yopq0bX/m+2h55yNrACmhBjRaRSn
N1yNgnEtHc5kIL7N8hwbWiKfQQFsxWpBWe2gKAJci9Ol1JeW2uD8oOIUn+hSJ4IKlpiv989X5vbI
JUkTdFSnRNYJJY6KJDSnyTsqnanwBTKDX0L8yHHXka4L9LBMDPNVUcIasfVVDifqL3PwsOrKTpuC
NI3RBjat0oJbnhxfka6svS6OMiNQf9nIjkCdxK4xLSI18449Au4jZOO2GEjF+ngXE1t/Klm8dib8
JFnocATkFAxkl+oar0EYLCnl40lMQ78KFtOkWvqsadfzaUOr3wiKTh0QiBw0B0kiWN/8LdhlKviD
/pfshgt1bhWpT3CShF32GyNINQYte94N6tfVjdhChpk3Ihwk0urwPFeM5CKHUjpO9PE/A5e6h2RR
PplFb+xAo+OXaBLLNCdD2FQMcUJMuaogspLqoI8O4NEI5sorVlxBbYuIZsqHISoaUaC+Q/Oh7MXH
UwbIRZI1dF67LxR4MElEfXsYYnHLW/ssG+AstbyB8h1/f9A5KD3+rYuOnbvDfvRhP+w8cORDSkTm
hNZqA2LSfdUqYfwBr6eoEt8qyJ13SP/XHVysg7ig8KCJHpmC7WlClwG04ge84ege0yf3fke4GwdR
bNOm7hRLutwvqmfiH00Ed4Cfgp5U0AKqI2OeSTh2iVFoNxStPEcrdffPHXNGFe4XIEt6r/eeZXJx
PDvDuguofVqJwsUIbWnpBO2zUM83uedn1ojGRjytz+GCt34jbAVuY0/kBgs39e6d8eTfdkQcmTmu
Dqb+qzGtlgweoFyga41z0ZUoA/Y5/kTbkExucUnWUnhazM0nkVfANfg/Yn1/VSakCqi9AEJe3JsH
tE4R0dCVjdbsjsl5vP70Px27AoOvK88vDs77ecO2VHmmyi5sStIEG6OqXuDq2XSOFFAwVHKSyL/E
INLakZ1Ba/Ffrb6QovYoGNMQlnjGAL6txjY2a5BzIEqyDXteY9/pLlwY/C1/pQOSatzjWDrb5GB8
JumBs22TKJyLQX7mKk+cYkhptQz5Q8cEDsLFYvoSIIkDbi+SWc8wvASF41M4W258bgOpO8ldM4SB
rjKWls9vwIjkz3ayO4JMnpTZXILFj8ICZUZ4vd/QNETvnAfy6HDu6MGAJGBx1YxKhorv3i1m5vJZ
3e2AtONGqqEe3znEeNFRVGM+f/dS7j6TSd3GM5Rir8IDizk5h2j4UzCZmGYGacwoYIrnumf9wq19
IlzpxGQmWr9WPF7lXOc40O1qDUQatct6CT8tk3O7SbnNB4pcT9+HPVPKx5bmtp5tewLgXtP1+9D7
KVMmpny1skiDZjTSuBqwh0W7htG6nLiWYoBPZa3hVnVRhYN/3+kE7ORe5QQ+1WprMGTun+b6idxD
o9ApOeDkfD61BiHMN2JQ9jt1ft10MOpmAfmZdmAHm/sSmKzvPefmCSh2WWbDbIjIy2L7/7bKQyhe
EjpFVgFt/JoV/wc+P+eKN6GhJ1Jm0OlpfVcTRUF/HZUJ1wpVyuL+d3OHoXCepbYr6Uelwed4BAtA
ot281UHEEFJIU8VGrHpYBrC7v22Bsfg3EQDNHT9gc66hdwCJG+R3/+wfhBN7QDHExtMRBxyUGpg4
YwsiH08EGoQljmm1RLU8hSJIGRaObK8Mwv1shHCqUM9pneQUczJqKzMDGuFJ8IWZrcHLrgMKpnhG
w8aoHtEzLDhBaaW3ceWGVnuFpKIyEgSd13+cvd++4UAcxFM0esybsC9bsR7JhYBRiLoZLPuAGTq7
2tKItINOrmSDqLMkIAmKGVpbjb1vAxd8dXUVCNNUzeaXol6DwgPSajN3BGB48MwI3dutU84XEyWG
NyBFRDDcI3yRDe6RrnhrNhXdC5nG7fY/bXOMBw2ckAe5UvaVXdc1HSP88DrFlJFBG3do0mqnSHnX
Sh7BB3oNDKA6eVvNVgGAW/HSLYXclwiHq20rd3vGnCu80z7QDQpTfiHxns9N7RpgMK43oYczDrhX
6RrAWtYa/5mv+6hPQP221/32IxuyrV/arSdTcgkPeK/ruvGIcP2+mgFXajn5aKAApUbnYbCP/7qk
wDC8hMdOtc4cTnqUH/CMrLaEnbUaNURr7hRWcRt1e4DHubKRYCKQlmoJaLJ/nSZgBupseOHRxGnJ
p9gPorJittKOc39e7kSnuLfXeYyXWz4XVY1aU7WvYX8t96VOe7bibr2v0FnbeT+Et4n3tTAdIYVE
J2x8NmZYi29xky6IBtQl+UaSaC18dOvTof/Pkj2ukMOWTrYCV32/ZoySdAi62n9G0R57H0Z92DO5
S6PZR32iJiC/Q5Qo8e6h74+BnPSk9ArA7/Mxst1mDafPzvCP6Yv7c5yJusTWGpvGSM+ye8Cvfpl4
8aAQcK86ySlMJU4GhDu0xwhCBwF8pzrwFQY/2N93S+NIZPJjWESiv1KxVpHHv/6XJwmsHItWk27i
2+vxWwJwnIiwFuzZr7hBi7T1bsSaCR2rtGscdekUbeGCxj1PNkmp2MZ1kd85Hg9Ulk+b/WLBA8m1
C4arKkwsKQmoKl+C8JUlYKjLW95F2j6MT6LQrltWyr6NIEqEklI0v+5OrtqjrXfPMe/dO56BLLWp
5+IvUFjSBtn724tQkWV3hwGTA8ZrxUgFf7Pxt2ZzUubYjpWp13j/FrYeADxf2KZODJhmSIg5+G54
ngseZxBMsD1L6+fmKeM4iozh/clnOgcJOIvHZQcXgiQeqeeBpJPVh19kRU6vLZbJgr+S0jbAx+P+
oFbQmeX1mYHP8z1KcaIMVC3PsZfXgwUB3wXpD/90WEQDboQ6GykqyzqSWCD9eJvEWJmd7gOItIv4
SpD6QLkEdWhhbJ+QWa5EbSWrWBrDdOqAYo3T5JwO2n9Ljd5VGC9D0+l4EFHotaSp1SxE6AKz1Ukk
gipQPMkqFhlnzYgYxuPcnL1eNntYti1rvoorHNRRkQMuWy1zztBFWwFu9ZQnCbSkaggarmK3pkHd
ZwrQ+W7XrpMHJ0ftnkj+ho3PhishvcF1P6X42AttbomT1xKO4l306zCBwhUIw8cZLUNqmM0XP30Z
Z/6780M2i3yHI73z7FzRch2o6uedKOgILt877Lw7NwI2/Zy+OmYQzLYyC/9/aBFop6i4GYBjNBBk
0BK+x6iqc8r1A4WXqAPP3OcgDfKC5Z9xlHzPOPDvzJqMBcQdUhCPEKnJaDU5b6U/tt8d2pSJjPxV
BPJ7OCrMBQ9U6y8R4kaSFwNfWOXi7LXnOhEH+BQNlRirB76ZTXvxpvw7UoQ3+DBJAjZf+HH6RrhM
LtU4XM1RDEFNz7oUtURe6onM2z5ZcyxR/pzzJCOqBLJu9LHrpY4jNecDZdABYMCCEbQIL7iUPDvH
kaTgOtpNL9Es3FEBnjArIZ28OOMQwiDGh9E8uI80IX89ce+mIE3j74NR61JNCbt+ZQDgIErcILIz
ILZGFKCowbb+RJoCjrcXjuGhoKvkAM/RQ1WTgJUd1OuVvVYIaZthvlrwzwM8t2Z33wkj933+p4xs
5+zeuHqiAGMfa7dddNwIhkFN/IkjqLjXniACR+2TZ/2twR5JMYpiJlfy3mYTAYwECqPrfeOwuGH5
uK+N5YhcorPuhjbHbxt0icAJPanCQ/rI07CKUPNXYEVqnLDG8BQ3mRct75xHm52MyEpgbinCEsCz
b0tShlcsjGTaxpktNwLkme/GXbs6THYb9CcIoLxVG+47XhVPMrEVfFl9a9wjcim6Ghv3fj59cXAy
vCm074Mgi3FkPdCRzXAPNOkCbTkXEeCWTwPy9DiRKqPpPlTqhU6YrR4mOO4It6rl6/2U+GtedHM/
gLDtfXG8/OPEieI6rX+y+XbTIul1Dy+GRw7VKQWaB4T5pdvm1evu6oPiHt6RP/imOJwQQAOWJdLP
YFXidma9RUqSg+YhpvRgpACcKLrYNnhOkltc/Ew2ORiD3rXGzahpFJBShFkOCXvZJCoVW5ZRQkUD
Q5PtFrBpD7EMDbTJFjyIugL1j312qMILuylq7rmgWGCGKxlhxz/foyRBA/+pYLU9LgQ9H+u8EASa
2vyCX2dELbKQTgvKLQlFWA5Gr/2YYvekrKi2iWsyjjUSVLzBVQCduFNuJvwACFK0KPqFgUxrU93x
x2+XNi9GlxLfHx8fSP1U0iQGZtWQh4COkJ+qRTTeEjQEEWFNjTr95nx/6ah1qfPtbwW94DxRuaoZ
tOmyy9D8vAz2c03FicP+tyXq61oQf+u3X8W6PQg4/pZpIsXijlY7biuC5m2yuurq70Ok/XEnJf1u
zwe5qhwVYHWgt5GgD6Y1BgF5l15WTrh/DOST/SDtJaWqUZTIGZcDfunwr1wfSiZo+Z0lPte2DXIo
jcvBxjvmb9p4h2PyZZLBXrfAarIdzCGTxmNLE8jfGUrOsRxOURyXyjMc+AUhrZx2nRFDZ1F/0xFV
wiKDyki6kf4b8Uz/YSLY2u1d4POWRcbFUAVpFA93vry2Xoc5u+XauXQ/reTJ8GgTkD2rwUzEZPwS
rhFb/r5noHlqeepz1CzNnWNYYoWPuN00niw6YCYADLvXD6jrl7Pu4JOzlTzc/WW5h3TNpcPB/ct3
/f+ix6bng+VmKj0bT0DRHK0FJzYBn15wl7noUNvIOBHkIVGZ8ErnPNyul6RWNFJrcfP0TrO91mHd
zgVmwQbCZGjEIvpGQzqEm9M0z9k4i7zI2vJlq6fIHdcmxMuNG3Oj7p77rJwJ2qPYXgCTvzxV9JQv
HrpEdN2qgNZhr9Uiv1dUx+OFDCx0U/bTbDngBRSW8XBznL38+6DWVSn93qQxjZObnkHXJRN5N21u
yBJ2vYQq8b+j/LULB7Ac4fcRfT5C1HcUYuwOxqQPP3AVy/A1+TKmA5NIpu/lZ1ayhmNDcLgC8s8U
aSi8ln0cX6W4zTrUwmeUG3hncWO1uAt3v99cAdq8eF5v2cHTJejfvFriFt/e9O0is61efIDodSie
zq/xLPmBCiZMVpS297K8wkrNAGIGqwoDcmjvAjIY2v2aeliryTwVgahC4GgS6yWEihgkfpp8hkaj
gK9sSMfyV41gfER3twNPAl6poJ7D6SUx+iTG8NvI3AQT4TMsllHHBmB9TUvVf3nEdmzl/yw6UtB/
JlIttcTOmVa7pLRUQGPS5YmrjJgw98H+OGPjtfxuZfQSqGIq75yn3ygvwQJMK17yoO71WvxLn4CW
UjAmzkJ8fmtJTqB4tUU5lOro4EAfIa7++rFatgmUvFZibZyvA2pAr6vqajtVTUQFXmK/R7UqwdeY
APP/Alg2tftFkbLi6rjpht5Vprvt31lZCXNBJE+tjzm6FblDwWL89lG+t2O/h2iT6Wyz5JAFo7gi
tNWLEtCqK4CJ7arbS1GyB0/vs+QtO1I4Ci9mS+reeoEhIXQCf0mTwFUuUhj99k1KW4TTmnCXyDa0
bkrscZA/jFfYSoFqnBRZtUx84M0aeJj+CGS+8hHi+xqN5A9kaQgqEEctVI6oyGhmH0rfsZo1rn5K
VK2KfpTaAgvsZmaOseRf74DlUYVrHy7JwN/qMGIidJe/jbSqLw4oMKpSZcTyvGLRX1/w6+XIsZoW
T22CQIy71iLL1snjnOZXltF7bV98m6wA//V0us7U/Gm0MgC/MvauE/0nO9lNoODHh19+Dvcvy9do
JP6q5ZuoGVb5ynP8GK+1pVH9nrzD0W4IEVKuYSlA1tMyDfwxwik+vHxc4JarhPXHESGqM+xgArzl
ASrwLifM5QnwhIrmhCJ1/HmeZucLc5d5SPd1kRNx/Llh2Lbe6fPLPklcAiddriw+RylVKsNNhEGW
bfQhs4bJA7Y1Z43eI7J3ZmB+Y8zzF1DVsVCx8WD8ZSfm2RsuGUt/UuF09FprZj78Fdx0wTGt0U5m
Jz+M5Wr1qAe/6pvoKaDN2zsrmjX0cSKi8wATW5GBDrUwcyKaCbEkMISXmZe20+OganRIsVanUPuk
CBzpUzT2YUo1ylm7q4wo2oWwszTVJLzTgg49GpkNqlCTIEgQUdO8U3PsQBb7VHSmn0XofyZydUL0
IjoCWeG2o40v7V/eimx0aX0e2TV2+m+L73JtiQ6DMV+4bQ3TrNoJWpL6xGEsMAI0T8w2q1b1lSf2
dylQfT67j0R7tI3MjJHVKKoJ4VMEwa+CuHUR/HKjf8egthpou03EukfFx2TSmBjEb3IX/Su9VUEc
Y3UbtyJ8dXSEL6eS0cleL8SlEJ4OP4MK9ffnlzxRApd0mbFxUJcKBv9CbAU8/981ATWfg5ZrL8RE
HfBPFGbQz9F/FeMfwahkcC7IE4JcmpBKyA6kP+oGIBgIS9C8SWw+VcM8nbU9bqm2X+oAYP9yxtR/
63II3uevcEFcZabyzRZxn+bha0A2Am22PMUhCUFaOxsul1+fMrc7qFdUOylpIVswwxNSQ9VHph8O
KC18oY0ZP3hNDpMEJYXj8Pk7+LUqY5/ZizX3Ju0APHB4gQNteV+EgSf516qaMPf5c2xZXbSIBVOP
tM8dVr+keaiChORNI76zqZBjPjwrhRJaMD/oz1d9ShFK+vAN8tMiiT8jY8MxHn2N9nLxMk80skI3
V6waL369eQ7FKBQzFSggaHdLb2XVQUPeQGegZTETHU+ta6WrLXdfmQs+Tlo05QS7KXrhtmyXZ9z9
qFtlLDnQLs72nmeF1e4mdV5oCWYSkW4tow5YxfDIOxj50znnGrW5YkWuPnqdO/XjL4KIR6VDln6Q
VQ2Hqmh0fMzdJ5rGEKx0tnpSZtF7ofUyTzVxfyS3qvgkeVITAuIwG9Q1hQHiNtrwzbOpc2BtByOc
9mggr6gzBRfk7fQgI1SgPxM8HA/HZHbi8HWXBq3dLrDBmGs5g6Xkk14Wx1uLjUNgNWsYzxZH0aYr
LFvRctAN+AjoLtiu7/EgDOZUc9Dvm/W//XBfeK/OuOsJbWtfK7TjAiz4i8rRHKWPLG/5hgRQE0Od
P+wQEmjCue17eO4VpkWHTUVuTMt3rmJKsYgpOFEl2+3BJbAgga52dYH6VLXshdSCKBjYAT8b08tO
EsaDKVzM2bWSYFYKhFuQINMWoATrZmrw4v6lqpZdlgrvjneDgrlgID7oDi40SlcO2XIp3jZXseik
wIcIHzz8fRdbsfoF175Wqj6xMMTXzMgPf0IcCVXrV11hT954rYVfsYfcOBVsEJmxnkVwyYZZiKVk
8i2FP1g4fbKs98TIyrwo272d3c+We23QBk2Z2rVhBwVb7mOOnjEV7Jiiia2h/2bX6ODPEJIhr2EW
qs8FlTBuYQnHMCZfQqQr+6qUFiYupW3Eq5DdGMSHqJZiGkNOBQ+Xl7Hjjo9ezOHFAJwDiJX1StKm
kKqPyvqzttkyBPfyJTKWaQo7C7Jjw3JgfE7yvk8Bagq2MFRJ0reHgfp0ivmCILskuOZp23gqtaM2
C9P7pdJ0DVKATk4abkAtlHvmj3agw1zVEM7IKUbsBwtzaRAbVnZngWobwn00Pe+1Mk0Rb3xjv7T1
itJmpJBc2+rdJIDc06seTwMbpqGCWkDQ4J1O9QjHOqNnMZ8wxybN8D3B5NhqVJ50PsdynFaZDGjC
Sr6OAwgmzeetDGmPHCzEBsyEKzIyD0JK2RMk7cNbsOhM+chhKrmjwHhaFF6yl1i6e4HElc3hEwxU
uqbT+VUp9ZiH0zM0Xx7y9d9MypA5a0zpGomObESuF7yBu2Ji98xC9wSjR9kd34y7fIOnwP+JNgEw
rVmPxJ6ldLU0gefUC55ft4L8bPDH7bwPJJbymrPVp80x1/s7/my33+RbrgM26Y9z6lsIRqFFGTq9
cuc4Q2FHNXGNDwlb4i+gqdZbZeqMTwMEmJHIsL1MgRfGQtzTPNmTNxIsogqZj+S3UYX7M22GrZ0u
QsPBc6LLgFLyilxx/VldXYjMYEnLQqFjvR+iL9k9u2Xzu3OfbolZJEI5NBCZJWlOPgE1ZxA+8zec
xft0wnFBMFtwSghJscTr8RRjCtS9icz3LkGop5+gUzeQ3vVtLZk/Wo6DmhI9G9Pp7ENMVKgff6Rv
V3IiJqOU3c3mAuTzO3EkcA5GPiTOgAfiC1FCuZzKXHSUdK0ungNQ0VIfkvWQN/TYyz8twQJgdTg6
FHMh5vw9hpyBH8nO4hMFl8WBdayJZtVCu8TKe5wmWQCsI2/WhuS65AH+JzZOvBOpEHsANkBQ6ffF
blSTv/brZTkDrxSvReFbxV2Lp63vUolUpYmXoFIkEpIDK5IBkT9L9EeRMxR3/RR9Uao48GcrLRXe
gxI55UUScacOH8+Om3H0LgebOskgdq735fDpVTk4M6i5aXAn0UN3gdzOCJlq9LiHaHoFK4vKNyjv
x1N5S5xMkao5P2Z6pyWJegYzSkkpqLcb7v6sIzMtpJEMv/Ah43cSxRTl+pa4c4oqtMSi8jhII/f9
Fq9DbEqTjBjPdzY/EbTZIaFp5NN4oQAdo6DIE4IFNHOCIiiHgXZQgpq01PSH7pndmOEdrRn4eZoa
I9k1BuAAEn5fCvkoM3x9Xgl2PgtJfppuoguIaiDyzFXpw9s/j3Rcxxb0JaAUMh37BVF1FPba0OnK
XFyBXeOpQayW6mbPnACMmxoJ1bc47cBNDBuVaSJT10Xo7TZvfzPN2creD2e009zVOazgoXeOJ9hf
vq+jevQl5b+XPrcA9tXCqM6Hv+J9KYYjAPseuNncVpGuSW72cWw0SH3s8+LhDw/qRuvwykLHo1Z+
xM6Jybre7Px2ml1cCcvBbAP98R0SmE6BPfZTjEz50E5rAPGPsrry4+kDW+JROl7m4P/KRpxqNTZ/
AtboloZtDOgI1vgatZVkv4wO3fKLq9RlMxb/nH2Tn+0/eCX4Y+GCBvlDpEnvZDQQ6O6SjxFRx15O
xP/MIPZphnzhPj56o1Al2reQlgSFJCD6VwLqazPTuQ85ioOj84C96VaQ5U1ddNmN4fv0xu7Y5Dh+
tSzLxUE73TNwEssX2eT/1LbH0t6HPL4XeJhse1IEIQSeBSrn5ssszitmasVAkPO7U4gIF7k3+lHs
cSc4ACbkvoGnI+uJo8WeyLzvFTxHD1sFX1iks0YoJqJDGJgdwDq0XSLB7XKQw8GoMhsMo9X83PIY
No5VgeKwdHCccfHRDI1gZH9KM5ufw+lmh9fIG1CjFWP//CBWtQ5vRUxGfYzaIw6CNao3Qomvpq3F
YyJR4DRICC5qatGPpapzaLC4xbxuOA2Em2blZRfYeEU/S2XYbPGzAZlnXproz5pvoN8AuY+dJwZL
TtX+WGlvfhDBIm3utoqgjTNwLIZcGj39XIxChU4k5zDSNN2igbMc/a8rNgkFdBbx9L8HCDhbtbMy
cjCTWs/4bQ0EQky3x8HVYeiwCCZb6FvyuVqnPJGsagcVkaI4t/e3aDuJnx9K2zklPg3/1s96B84e
XTc/wvmBkYFZ6wXVU4Wlvni/9ZsXJ5tXNOH6opJNjCXa/+lGiP6T+GWpVDaJdhKJO8Xu0mrCcYfQ
vJP8HbWzeUB30oCVYU+azKvEhIKrd7tgY/foesJI94C+bnlb/sVcYgmBsBnr55rLiUqM8Kfx9GJ0
U6+f1++4g4QBEmnTK8I5QyJpnFMxMiXAmj6Bb1iTPS/dzUWmrcD7a2+c+n85a8vP28FkWchJqAH9
TVtY9n9cJszWhV9xLvjBlp9I4DzKBopWrYIVNtp48isO21s4UCkE/aC8mUvr39AtbRz7tSV1leXC
0z+LQiqey/3CLBGCxrRbSfVkGdGnDuCvQ2DPNsiuQPXgLfWqUP+0Z4Tg1sDcsy1n/aoM7PKsu/nq
hhFjdqRZ9xG5FPW4UODTk9X+WWv4TzOnOsMn0CpJ9VzsKoof0L9/y5+EHgvLBjgDdbDLW4L/nha7
gtMawQ2Gy76VLd7EtJvwJPex34bj8ZEYckj9vWjAE36k5bBt7qRffEZc5P9f/fse/BgV0xpo7fqb
KDHLamPE2gIZ/GLtrZ16Ffaek7E2gtYhB4FnT0tb5sveZYNnh8b9aYdK+ScZ5eB0ckSHdalMq2AK
ywsw3n1lknqB67w8Rlx7j/sQQdnRSjseiGxBVdc8DSpFrMwxpBTg36V8zrhS5OjJGK+0P/L+MlLk
8EQfjgkTWBDX2VcGX1ShZptooED+qYaDxYiEAg6sqG187ZGXLRWLik7A8DKUkeqFkIYGo/RpFQZb
zZoKKAHkn7/xcbgSoNRmzm0JnQycECN/4Cky3xI8WLUaarKz2+I9HaoWq+DrFg4ME56FYNv6tKWN
NM6l+HdVyt6ReTVCyHkXguZ3j95dFVMUb16gwgVYFu9lXT+Ox6/X28GxKYTHyiIoLNSNCuYehZUb
9P7uFdJS9fSY+AZTMd7SoHGaMCOdR34LSycWspbMTUu/7H9chWfrg6px+hhYi+tuWeLNyYxTcEzG
gZ6HTHNp97sr+5Gz9H4PsRPGi9e4hrzvHk6Okya8DiB4cWCvwLEgmuKTPZHFWsJgQDJ7g77oqI8u
OGG5LD61MXZ9uJl9lTg6vt+MSo28rk372yEXB1WyUj1iVMVkg1sKo7+OMWd2biJnx3wJ5xFlRo6S
LatZnVb5EkpVDZSGeJe3aRA8py/pWy+hH3x7uZT1j2qbBXOsopEGopqJgHvU73STAHOX86+h59WJ
jRRFBMV/Lx/aIRuf0XTpd3v0lJ52uEQ17YKj7g0qfOMzKGVqxBiKOYeh325JRZGKzwk94QwLji5G
Na13CspWV1YlZd35OiwXuHh3l25C9ZMZkh5coe85+VgFpkAZ+GGeywPSWqDCRnBd3glEHGxy5vvA
tjZcAaUB2YMgTKoffVyY6qCjSLhy1TWh5g7jOuOM10q8L7c2UnS8uudNmceIjVG6EhT/uSTz4uxZ
wirivdpYOfAwAGlXr8QKHaqztLIZxJcF/FW9z1CFUGtuAYKzF9FIygw0IDbTkXShgAC/vuoNZcRl
GPx5bCHRiNDicTdS0mjdUV/Ep/t2a05NDlNco8Lu+yez/NEE+onhYc+e92uV0xCphe1SIdF046vM
i0eyZKxwv0OuNdCT8cPvxr6x5H32KROXY9LNsIHlZgac5fe9PISrRX1TX5+k+ZZow5XPLSSAjrW8
tAq7iLDLasEMRm3zZlMLcetG9E9/Jbt5lm/bcQpylr+PVOVQaEoqWErFz0vrnThLTdR0BGOCDOAG
5qPsMDzIuTdNpMBPmzF1pqWT02Jh0rOfE8WXE6xaoeVnmmuUmfgKUVzXWXKggR/agALqK9Rl7vVY
KjnTIEpymPHlIHC19q3WsA5j1kZyFTxuesJ+MXSL13emjOXd5ouRTxgK4pHNuc0wW6BwAZ22ueEB
BZtc39+V6ACO8yo6KEixH9uB9WpL/mtGt4hSgUONpy2rm8N+puz0if9AgxDjFJ0cPNHrckGljQcD
Ferddi0/xHBNxOgsnz+ibSoH1AyfbfBe6c9DAa0ZNcKx9LlGBfGDbaTIhQOGfChRTLBXrQy3J3Sm
SmMoPsExID5tHtQ6K4g59xOWJpxYafBxtA1TK+32r6OQt8z7RFHcwdUn58Da5W21oIEwHq8xMzZB
ztj7fYhlMx7qPeJAbhM8ljzdM0eEo+hSxT+eIIgSTPfcYVeqGe16GjtZKFktjnllj23StgSd+jo/
YbrQ1xKKvrzZmuVWGN8rHeyaFOEwQYf937Nrj5VirntsRX1PrUhYcrmjdbq2zBi1okUjv9/hFoz2
c9a30h68du+qKqGsCazRFf6p95Sq+HEPX6yUiZ3AV3dMelIeIzGEhHDvuhNs+fZmAsySlX/GNsn/
MjGXDl0Js2TKcYkYuHmxnTFIXk0J7aSwwkzcJTsZWTzlocQoJX5gyG6gjBPvH5of787D+fSH71bI
PrmN8tzkuzbLCcAVLTSzD79+nGWibB9yfZdpL0pBdG0QdnyDG2ZNvC7LOb8Ay/8NXCCfuwkxlP5x
UJ3A2RNxKGBhbxcPWg7FxtYUvwY2SyEinNwVYdRxhv7EwdlOl31QWMv7eCZ6lAJ7A3y86vDB2icJ
Mb3xZbJpNQhNWiH+Vlb/cuwuGoUdvdzIjKCbtmoME8ocGY5jNFw98xVPP1+A5rY39hRM9/PUY4h/
/542cd+cWTX1Xa4E69ACRpVSJemnAOL9GdX6N3acxYwK8Nylb6I5o0k7wIQJoxgJ2hxFr7R0/ifc
mY4dK+HUR3Z2bPPQmi8ZZ7U7Ajmno83MkhkNxPax2Boq6Vh9WSaqa1ugIb/NUJpLhT34gFHrIreD
gDtg0iu6d5HWt6Z3fVy8y8BbheTiNErYIReOTCrQAe3K/eE6IitGDjP3RE71B0qzdGENp07K/FDA
uNCyswRK88Z7dkiAxqE8hqLu9Y3e0cApLv5I+Zz4yLg6cSLS+T6lQeER9sOh6OWcwUINcaODrReI
WBusCboPNE+iuCI4XgfUbmgG88V8yVR5jCVzhhjUYEJNXT7nzIrITl3FVxBs24s4W8X38kQknGqf
84c2tOiSSQtLFYh9Yd+aRPf+11BsQHXR261o/Ehclxc0ywqgKqg31AYhnTuaZW8INABAUEWzVBZm
QUjSQ6JDUKcv7FoHPmnSpPQuqXuekrcOyUOHtE2aXrsgya8ohWn8z5p1G3eelGCqRYO62lO0ZnZx
WyiOlmFReQmrUEImiHNHBJ3hPteRJrP+z61/BcpR+OIf68I2v0d0TjBNbua1T+dil7GJQUEzSRdi
QrrPwL+ywqD4QaPDvPCGb1AF51Gv4Ozo5ZGgeKs1Epw5YpRdKuSgiPUd5WyooBCpBGedLBCoBPEF
MdVzWVn3UGjMXHJUFTLotwYBUI3bHS3tx//jFxBvAHcnQpDQBM41n9KMgLbmVn3RUxuwMgxHaWTw
jRMtr8qWnbQYkB2imJfPcWnalVwIfJ3EMH/4ZpubedbXpcOq4bTjuIkPm7Hg7mgOwtkM1vwtl7eT
dSqiE3Ow/RsVPSwySpVmMj/CHEG/BEgyEtLq7KeTMFavIA6R0KUu3C/CabL3p6E44dCmMvg9LXfy
6TioMVDKkpzbK0k6EUkLPjD/s7PlLDBVXW8dglRKcRZmlDJ8Bc36cLGTDllMFv8Ei9H1+3i87HtY
feOCQmnNzYn8hj6yd90iaBOIaECC9UmUTyuAX11l3VU8swW6PLk5V+Ch0Jc1zx2X580kMDtOUm6q
k/WqMTfMZ0WcfQoKXzxTEHcl1RaSnBlKA4SXPkdxBbJoUuzjgwTYn6qihFTMsceQinEviKURv/4l
q/CTuijwlu4G1duahEUERSbcaFodtfCxUrCNdslYMSpDjx5IWAiovE8ffbNOgQbOBnaMAs4BkjWD
o0/S0agcq81OYcFd+wTNB72680TwiFz2ZIs8sYkvuJAfzohCfRKJKpHdlghiQLE9kzj/sv8OuT1s
AYNCdSCcDTNIDdmb/9ikLq4wgzCGFjFArqxtynKJKfSzaHz65GSbaQrHxLvpu5MIJRaLEYYyUJ2F
rr1zQw65fgd2PjwMJU/dHPi0JUWE22/vaL1ShCChbIDXnJoJCD+NreMBMP2E4x2M3NnS9+iFjLn0
uAU6nFDEAhAoa34Tnu7ypE/3Sxt2MLudIJYuZ7Qp1rU9DtfKicdc39mxsa+KKBYDKAQqC97XWsYl
yxsKliegqtx2LilBh79fbSgboDl+hK2u9EFIgdyRQWMTsdOnUbJdagT3LMs7o4MRun0ZSTnZyIun
+ZF5R1Gf7WEKEt/yIqFs8wE99I6g9cHMEOlf9U9NOmmAkjW0RzIZEIJpCWMz5o4Q48UiXx4SIODI
67agfyiiD78gbocIOf6Ir4yooHnXMtMWsZ4nIK2p4NvK7O553/h7xlc83z0iFFl6I7MAa5jaDoC2
AFUXH2duv0zhtw1TPQJc3xJZqjaEgU3z+1/XS29cGI25WgIMPa9+oPHgnB97QkPH4qlOiAFgNtql
jawsxxQOmCMW9zZPMxTmvLpdXQfeswq1QEVC3wvzVm83o1ndpT6aBf/tqByQNVIV26v0cj0vUako
tTcZDc9iJCEjA3GQy5guaCi8jwsZCVvKXYmHthgG2T1C6JGUZ7AD63Xhep4kZl+HmifJ+GHLbjz0
JLxVZzUkakm6Wgjzdor4hh/j+XuHSi4YXpCSPlIp8V2vf6jyEKEZWSFgNdUntArwDb/zr5vpG2Yd
GVffhVj/FpnRyZQ6A2C+xDjo/8LrZfnD0qIPn+H1hcAz6FTZearedGm/t+LbPKmbbRX+N/XRaRA3
xh9PY+GYICdMt8O1QtdFfjAtaokELGLrjTgc1mHGokipREE80HJ0RhO0sUGqiqBbfokAtHUawhML
Md+2WHIUXZGkqBRwfdj5RdyKzUSs7kxEPTZySUoZYufSrwrSc62QIjEwF4S1sjSjfIk8e1fJEvj1
WFlU4C9NoNLGCP8A5vAL/lSA2yZc9aj6t43q0v2PcFCxTYyxRdFdIp5Mx9Ccf9tiyIVLneQHv4xV
T5KJK3m/N3EZFM1B6Ik+t5kfSfpDPiCDSvvF+mVXBPzavkzRKnUeNSlpJljH8L2rNLb42mj2g+s/
y8Oyl0f233AAGpzJSlxVbGb3s5bZ/b54Keiy3cu0S1vjCeTdsJCF9rb61V+hKNZqHvPC0NLp2FS5
OrQJOHWnn+RnY2iRsm24F3mQICtnWj2Z42yS/CQmLVBkrAO7Hx90kXgjBdvzkSK1OzMtjnz3V6JA
SlBcxUCehdaiXMKmfDswGwttay3Erm0R+USNch+/vlAECK7OW6f8r5PcKGNpGkjYEHkJMxgRvQn+
DFHsxLSb1m5wb6YhlCXxgRXJuWcimgh1UTxxV51PGed5ccHbANQnV2pyMHTqE0LrI3UM9MlVmfGI
hwTCCvqhuBzBIt3S1BR+skpsyQyOxBLa9aaVDbRTIZcGmx1DQBC2l6m6fJgrsCCyZFGwEQO/XFMi
zQbg873ESG5+g9G3c6IM3kcqV6NZwl1U51U04kTwmCPBWqOuhlel1sFDNViW6lIFmx1fdrZZDe2J
edrr+G1/w9Pgstg2mINVudsZ/eoC6TBXtZ3OaRwNNbxm5H6FAadyhmV9yDlQT+CaCN/idVBLhKh0
gxt8AhQB0PQpIJwmtk4pMKxBNF9s2LZVpDTkYB5jhb2Zy1RX27mXP5wiuoxjrGbOojLJeys3e8wT
6YCbqUFG6SW6gxIeAJQ0KWz6gj+r+xVYwIn3ZSorOLsm4pjIKJfUtv6bQfJsDEO47tgk2ZCgmBTt
D9YYTxC79k38m5eBwoVwCAK5cy24NbZ46DBZvs+66vO78Rg/9SpksfztdMlwgpHFVk3WcITsY4tC
9WoGkpSNSxltrF7dDeeFT8Ii8kRhkZbCv+x6Qb4CdiS7tS1exP5RQOC9Ps28wUj+O/G/cMX2TUkp
aRBz2GAtgqs3H1CogpVKlVg2u1XBGlvRogOf45FUbiKlonXycasxCIAtUK0aOGhzf3XaF/Y8UiF+
SlfPdhrgjz4BV6I1z9QO2fnAk9rrxx07f5YvvRjnWiJLlzgIrb9zFgC7ytiGAlSsYloKiVsaPgdo
BD7O7Kj5Vy6UDSdwm4U+DI3Fa6rbnvfCpn/j74gKan/lgeLx1dNG4g7Gzi0kWMLLd4EIe2y7iBGa
iXmYNbS2mxpYY/mTap2uZQWBPDU9+gdm1aMpW0vRqgjyzG03EkOVVekno+ExdMsmmueXmMIMVkvn
2vD9r6+iqAOmfz/0EOcs+F/H2bEcKOSQNeSlba839wd2v9tpKxKbqMKfVZafusmGH/lz+N9eo/FN
GMsOqU7/Yf8BKBAbVwLPUMJjmIATj3RBzjKn2NhSjKwLAZeBqZ+dNV/ueQMTr3CHL15ob1SB/6BX
MbSnn2DhuwKOoe+x4wNw8T4t7Sjaj3+XC1vuFhB8GwIPKaT7FpYEAG1kEgso+BNIb+XCoZP9mqwW
3WHZ0J74a453Qs9zuwwbKbNzsHrqfo5KI+VUzXP0ANJpavG4RpeRZXiilyb+K7djxOjdTU87l0SG
6/pVopI4ZmEeJ1a7oNJTwQLuJ6eAUd6D4zyz7C/d7sk0juQ1yua3ZvETUdTFTwa61WZnJq/FlS4u
2ZmlkXyelJsWhtYEb4t3PkGkhKO3mriI7Yv4L1qZilow3dKigE7QcX1MKDM1bL21zX81jJ47uxIt
AXBNeXB0o4iFYEfqur7UwDdCz20KC6R5AvdI1SHOheAtVFm2E51ugmefEiORJyZIYYd2oYzeOjWo
Y0hwh9UmNDZI2TmiV+jomlYK+B8/R3RvID/acEhFFk3CJwDECq8lDmw3ik6Hz1nP8TS9M3ME3YKM
4Nd31qkPBeI0Lsk+IaiMGIybtnid68UzwJpzHKalaX5FYw32RN8MDU7pVihArx+yZGNsyXZkm7Mq
Oo96sNGHjqzrNYQsBtfRAd/cglg9rTXyuX1VsLLuee4BD+6o3n4YXfJcx1iLHWtypSvpvQApR1Le
sdq905n5eBkJDwYero7nSOQfIdCPlJTIzGXCdDf5rc9VEDJ2CzRAIafupvRwY2jMxf480v+hzajY
yoRIxcKQEve5/n1SFUwZZE98U6r2ZErkIiceUCAdmCbMgE1AjPuKZsApFRAm8m1AdxY6jfmSKZSS
VetTsoHkZ9/GKPcyXC7QzLaAj8UiDGWslK2DK5Fq8hIgvuLPzrfMvUsQI80XP+6xHfADWeCKeugJ
qwB+cQP+S59KjVk1lW5NRKBKksMsNM3hzFdSV6lPAtyazccn3gsySwbS9a+96UId3fVnM5bmiQuA
KiidXkbL62QBLvvO/FPyoCgjBAKxG+qoa7iLcYJ/0vDB1/Nd4wJHR0fFAZNJD7k826tdkGnbgQWQ
LMN/8VwxFTZzpv+JN7Ez+2DCT3aR3Vt1Qv+IB24wsNsJUrJPoygTTiEFVr7hOXYazt7n9huzFvg0
ZesvBYQcdxmfLkjc5vclDUc9aAGf3v14gXFZOzJj4YmOSDqH9VZ/5spSD5SiJfFl7IRk7eKZAGUs
3VV7k+tjTj43M5R0y3l5pE4J23wEQkj55IELGYQIqFE53xAuCITvhdcvEjShFt5lMwqti7XiE+E/
Z305n4D5TRbGTTNit1HB4IxjTOfFq9c5LXK01Cs8d76CLdWnCTUgvYCN8qZUpOsI49MdKkCULm0h
K8uksIzKxsE9yHzu+JyVaQIEmpHKctJ79JqOAaIMk1ORt/PwuZ+7jRbO1Uag/vcu1XuPwRt+oPKP
9pukQSYXtjSHrpV5+qXr1o6zfSIDHVHOV0iGRf0TVtdNGHWXpFK7WUAloJtwYAqzhK1KDCQ3efOd
aR9YeB+ZFrdogHVeiaUsLCCvfRUinLGhA7IH6/hj7XjNR7LWM4GBxiH99zOhMRJIqn0UtWDKN+6k
8Hd5aAVaYfV7jUwDRFcRgvZsErRbCsFZzp3q4sPPUajl4IgRF0m1HB+tlIg36gkyp1fprwnIEobn
7mVBLRCpfOO4QPk/n++li7Wk6qqD0jZkq07MxLvDcTUsjHjVUyywfrXHBHMwuQzidxhKSmtycMQd
zcg5MKXYDLGucL6wm6lWG/r8bqw7lAwC0kv/8V7ctbDDT5jAO2eYFIu6+2ptWcPHsmQxwCWXtwT1
FKUgIY8hH9+Wrzk/bYibYhP0B0TQNO6CDDqsbVA+zeJxhi7rGSX34b+PCVIthCKSWztV3XXv/h/d
yIKl2EL52pZjy60gQqFnuT4pir2IVji/w7rLkMfKsc5TnF7KYQEFklz8Ap+BtMoMp8X6v9U0OKj0
WzQR/V47L97GyW6L+urZJ2P3elCvgQ7P2JAvVGutGhtVVZUhLvNIllvwd34y9ngD/KrDYbsLzI6j
xI20dect2jGUMc217v+VSkCpakGEm+q1W5SWvcnUiT1+n+2FkiRzXp5pHovek1u6pHX5n+EXBXzh
y+nh67KareduvrS4wYL/Ld7KtDWIVqugIUtPkQlGou5wygSvBd/px6mP2qLc5/4NVwPcjgK1If6A
I6ajoiWNb4zMAECFqgJZB/Rc8aJc06QZpFJ+K1oDFLVajyXDAmTIorAw2YetlDtrGUiTFqiMJHc1
t5Zc4A6gn/5kUrLen/jUENaAyNAMWbxNp2qbABIKPJqefqLoiY0lLM8YV99az1zN1KxTaaa/4ZEf
dNawb67ClKvxfU2PK5HpYROIqT2HxNnZuelItG/XKxXAP4L7y7dW9HW+3ru7aNwOKtwfa6pCuuFf
QfINv2e07DgDHzUphNVjsnnhCZCdIz+vp+l9PokDHFINDLCEMvo5e/UfJ7RgfBykA3Q5zYiW6kZm
I127qx9mfy+ELMxcnywkgRnp5NQCFRJH/6lfyCBnUiqcWGrR/tqjoQKKweyIwqRFPZosXED8UvH9
RMdf48O28l41AHzXkBXkfsc+bEqG0RNO/nCfDmjoTLUEvrlMRHOjQ1ks1T59eIduPSWI59OBqAcD
DXDNrzQv4wx5rK6kGfFiVOBEYXSxncjSY6Sl0Q4XV7IRn3yzqyWo5BaWi7+s0GEhl1tR0JVFFQ9B
2Qfm5InL3iDfYjLkC7je1lSJxxmC07MMYLiaMkIIxFUhSweKKe83eMmTTr1LnhbhJEAUYbyss7hq
6w/aNdyANuVDb9v4wAkQE7cZC3G7CxlpR7c2gQz9qQ0rbCdKVyYILjJ8wKZrnN/qi+EBBS0PDnKI
J5fx4bZ+4F4um958hDn6vBofPYQbrsdwq7NDSF+dDp4YlkaN7mxZ0pmhhpSXXsweh8fdsw2Dv58P
ieJjIru6xej++5FuCYdIrij+tSKAYm0rsS8bpXUADwLH5Nb9zN18MQjgkhAtditY2qa21n/p6oB7
yLc6gugqJRmzTXOQvA6Jlb3Sd4nJTaXagyHTYZ2LunLD9rA1Ne4TyB7uNLkZ+UprP8PFRYGzEw+8
fZA3MMrm4fEQbiMVe61/81LKJrN/7ZTpkn+pncNQkY7fs2ltDtiCaBivNmv5G3ivCqfyGLN/r4ze
nYGmCvgiy79/HqHf1jIOrq4WYkemqoUAHmxdal1nRDbkjEYblrmfL1fg/hB41wK83tpLgHbZY8gC
jc7PMrEGRZPDZ2Jf59EiODbJDeSYgKhq0E0RFHGOLxQ4u51qssFVpj/xT5AoQ7S1KUGk79hg1Fvo
DKyr5Cjv7eJpNj+pVWo2O2GpblIIcbNIHNFE5XNMWbgceNT/lEbuobihPuKTmAPrSjsh/+c7K6IJ
gnkF1/6b+JMBcJRWnQz3pE+K9AUEbj9+7ys0bCn+R33arBTi6H6a5a4xzgD+K8xO2N+mxQlvuRGf
UPG5gz8MmTAgDEA9ll6rjYG5Aj1bSTKEMZ1w+h+XS5XrwJ1roFsPdMQvSVFwvPLZ/5xEE+7JiW0/
WUUfv7kaU+xwqS2kmnX+PiT1DRu3Ryj/5NEkpGsit4fo+s/ho4fBbprgB6LX15STDOV9Rjin8P8v
1nA0TDy8/JWXD8nvRUMbQO6oVeeOeuf3RvF/MsobJfjS1XcJsX71yH3lboegmKepwa/+8in+wqQO
U3qXOnhdppCIu/X+p1GSXu5YydPfIjgb9Xg7TbBEvptupB7XT8n7DjifFOFvfgx7Rg4vVOzy7+X3
BQb/sJ1Sd2qtTvjAyMOEh4RuA/HjpXeKCKxfQsCuy0S7qkahVjbElzcWQ0bvOZ32OBBHGbn+VCwg
7peztvv+jtpScHkbZ/QtbWXV/HyK5LkXWBOtswxPEUEDUpHWkr2EzyNP2p1+8dP3bQQR8O4pEMrH
+/A4BMM+8Poc+WG65kpy0lkguAVHM7YWXABj66vh3d5lRCYWSy9GcnBQYOMPt33goEQwSHDEitFc
ohf6zDytrQEh3i60jmXdvXODcc7w/tkDQN0SW+ddOIAhhl2meGb3lQgEbU+CH0vz43i5jQHjKWYG
XNp7KpWbg1+S0umBLYiadp0sqDznaWA9X4p+Pm33uroRwm0I/in+qXmrQsKwY5HDoWHGVUT6q6d4
RtoEkies3yU0YEl25QP/O5RNkPHCCIZcSSGnbzr1Ln+zdrtFXfQ2RZ0cjTkG25qtrYfTBb4+FGwj
ytqv2Htg00rGCF9WJoo3Nbtrk4pG3UukPnmZikLDjKKOfhPNRU3KLbkzcb5SMZPrNfDZRMsfwDnI
4/3/duLz9nDyaIAaFXj67rEGjh5OHi9iN8OJlntPEV6rUnce38GK58BzJp7LIIBNCYe/7mPFJp5p
mCwAwFcAnDJ/VbBOQVaZA0AvmkrcpdEVO4LmsQICO4d3Pp0SGp+5SGBPhnNQhS3ToHOxiQXiXiSM
2u3NkBAavMdVN+quDMDlvI5xQ8YK4Wej7BaPq+aBUrYYYmkm+bKrYubZ5JgAy8lRGnKalE0WL4bY
KDvSncv6FQdy2O2sgxFFjbj6L2BJUq3A/wL1ZIBEg6/MXi54+/FxVpttZBcTn9kxBwzvsQvjgop/
u8FPV3QuZxUDqjV2Dr8GWu4HmqyHZ0U4C4G6zx+wtBuDssSbPgMzK0h6R2z+Iz8yXuRxrtPiEsrG
YD3zR7j2remX4T+I3sT3IbmppmFSkTSwCkxJQG5YmJOO2mdPZ7PYbxA054IcQgpGbD21d53zvgKX
9dUx+IRfAxQw9A3KA8mme8QTChyLqUqm8Z+voxDUUcdmYwIIE5GU1ou8Zeb5N6z4Pz7HvZu3aczx
j/7WFZkYRYvM5zxcE/ufPr+BBBBKIDHFmEmdHScYFRNaW8eZhfQe6qEBw30lpXzFDFXl730JGrYu
8kG2yFYWXk/tK+xFY+pAqhBZnfgrGr3ITaih4OHyXHvALH/fzR0e46ZZBgdjwYgQB/i2DAdlQJk1
VULH//gtRT3WUxv52kRk7BHKpZqbLRbKQuieRo9leB/d6WgBEr0C7L2T4b6TR7uTpRtdy0Da9FZj
dOqzRyuAuj+o13Q3qJ0MY1P1d8s6v0e0EdoQfKObpoMC294MVMYMMMC5o6RbgFgwsbTmXJhZy/cW
6dkgU4S/DDHvx9hDZwxGpv5v8eSQWJJrVNNYkOrq6or/GidDN0ztPA/gVfzPUnuARhEgEa5yx6Ie
PX3l7+lQLsiLt4MLdxBdjoNKPEin/jMMR14bCmSW8ZZihGDRXO5yoRh17i8ej9it7F/8w6quhwsB
oXJCXm9PlFIpZKHxhUgu2U38OvvMmB/yY+IfJgKFD4HKRIgjMwVjpsei9akcFTVyiEHmywYYdTbM
YrZ6Bo5C+oOfR5KitfxUJK8aYJGrSRmQC/4EbQ4CH8IoXb+Ws50c0D/XgL31wcHmg1IFyD4Y9cuV
sIhcD9sWwSqB3uWGQ2Ix0y0fj5XsbuiPg8JhNTA5Pf5If2H5zLWaqXCQ4vG7sL7f4Zf37z+/ahSn
xIYG9wTgjCLLDe8ZsVH6lwUK2eRwZOZ0GcD8nov17b+4CIrJ+QxxD4t2nciedOn0CCxIwMGj4faY
YCKHrvXMFLsn7xnR8noQbQ1XJ70nUGaDwtsAPePTf9+2twPzOd/xT72nesot1YEfLX5FtKJX5vCa
xn6p9/PY1D/SO6wX45aA7jkPDF2XDineWr5VRwrMQ7fLW3KWc1mD8R0Lb6iWKcLZlzm3XQU+P9Bk
FqioVFRAJgOigr5OuSFbbtFw4W29dMNe0q0ALZLFHutRpoHWV2cVNJU2Akp3nKrnarfQnmZS2ZyI
cSp6bf5Ty7OHcQNDwDZwtjjsRBuEcqPN7Wo/y747HSy7XijKG5mvL81eo9MrcwW4AUaPgTTVVyDA
Z6yII8ifpALIgDMSeMbRISnFVh8w0Yv2mxRs7QZLrcNc/jmZcrfRJhMHhvEsniganwja5OxrVRbO
HLXPYdyR6yz2ERDJh8PSYFDW2CbYZlEMAY6/js35iLUkVCM3Y2pfyzuXYo+WBoEcVEsBnUXI3y2n
8YIMofSKAOMVZYB/WfnyzATKl69F+4vbfL/zJxYa1XD8F/G+HfQ7A1rcyzhhqqU8Wgw24IV+rA/u
c7GnwbZGiLqfH5tlGilUyB6/bQUYHB/jCjmTAr2HYZmiZvk/gTfyrQkNczYFVUUB4OIw8ia0uRJi
opqoxCrRBKets6T5/eMCsh8cB/M+2Zj05LVhgaaxTscpcYJcKc+S4fsALVMd5oeXVZ9O99IhrNFX
vf5E2E8ffvy3YlUfutPN21zDuzV/Di3zzzIYt/lyRt2kUJZ7ZTaNrdKzMSjjZF6hyvJqU4PTkw8L
uzWXo+onDeLjlDfqhWoWXnj16J75KWAAKuD7gQdK4MMjNi7e+BoTv9qRA0X4EnPQIXBh7s66K3N9
9iq2MAAe0mQa9FGnsngJ0TBUnlo9qKvf1ZqHzdFTxhGf/Wpa0GkrTuyCg1bsDj8iPS4OqTlO/m5G
KaHGe/Hq0n0OxOu0gdM27/JubWRi0DR8gGAQbn6wuJFeThmX6bWnDlRytYvOry139yIgYIcEM92N
zAHa0PTtAKCqVqkuJhs3ZYHVejHbK+m3ZQvMCkDtufYnLhJzPorJFTAVtfqndYmel0axtPmrnXVB
Im4kqv8s3glisyxzlLMyV5c5nGOcW00gHqEk9JE5bsPArevGbaChKL2YluitRbUcU6+7208EpCnm
uUM+/rKY36TfM2xlk9YiMxicQgKtZTbY5ssULphIXee14mx+VB1ZmvsubrPuMjh1Rf9QJWP/nMtQ
+6dZ3yxBYdEKgE4YYmRQ/ORbvnXjI45ZJzexKWwWEWiktRpZasfXff6NHkBKIShs/96JOEelef/q
8xJ7T7LIv5pN/WxovxzPQsALADQoYFv/Hw2n4RqM3aqRVuQpjNl/7usdhapcvCDslL4C7jQb+8a/
sctOqSd2iLabAeo6RMQbNc5q2mE3s82PfMXGg23SY/H7tHOFEEg28hg2TYFDusHCqTm3MzHA12t9
wEFiHln4qSLHA/mMYdyOqKTeAsIYnCDzl7KghuzAkDAm73Kkb2hBQzYzrHC6qgCsdqizNfb9X3E7
wnm509rYOtY/HKR/HElIdUH7gUQCHmg0lZS7bEQ1Cv7Icq9g/2C/IlQenTI1x8OYPqr+ftMY9hk2
izUXu2jtUrmOuF5KsBN7JQMhEz1psecaZNtBSM1NoKX3MGp6gp0gj+KGzZEEpBBW3fzUbWuRRtB4
f7Iw+Pzrid62ewnukbAXJ9+hGiDo3ReoGZsugDugVkl1K295sFRFB7LWYDut2MObybDt48p3HJQa
KphXhgjJ6xzLqph6SiskftsJb5KqOtoa7YguZxXEWpfvPLy32fwh2E0Dqdy0mDK3tBYuwGQSZSSx
+U16+kx69qh5ZoPqGWB4+/+OKKpemTSFJodfgCckwdoVa9Yp5L5nyvl33HbkDQjgtLTLNFyc4AsL
Kf74T5mFQw1/muwUm2uEdUuyYpdWTGBu1KvX49nGMep3ujol7Afy/gDvPcq37V30U6uiX5tInzZ8
dihPdRvt5957p+xtHiPqENfzl+lcpJ+A5bvaL0nZOxceKn+FjyVBv3xCqtDi+T9hdQxKUvYmpXVH
ZUenZwnZpa3tRU8a29nCtKmaAtNIloeHKX2TOcgHk7FlQ/4261Kt+Ygsuf7ZOxq9BM6Hc+EMLnn5
m9a4/InjXjdGnY4Chus99GDEAzutkK/UPK3Y8Nicq/ckPFvDO+VdctQDedyvKop3+TacB7SkgaXC
UdIVjwl/46PcTVodcJ59TxXbMHoJlvislq3+emXw4zQX/PLtet/5h5uCCGV6/zkbrwOhzjw8DxJh
/dJGqwZKYvn2MJ/KOJw34f5J8FNSzGU8GLGAiaAp8GYaNmrx5SXvGgCrpNQDYt/oWMmaLThW2daN
3k5zUQ/w9+VeInNVZOfcTGuAgyPSszpE24cZ/VaMbUxJbvTSujcXv/y5aG5I4wObSUT9xXDC60M6
pLQs4od/ehWPjYdEb2zLT4XkV80Elfc1akhoi8PP9ejhR1XvZ95mrYjLs9tqF3n+Iorjq+fz8fGL
DxG0ekag0dBtMrBlTXtwxJwBvg8+brARj0y0LV2F8+g/eFbAy6k+beacI40hgTQ0NmwZMtMrYLoj
AwjkhixpDN6/8fudE7BMJLk2dQLfc93Lb2N64Bb53KHXRqWkAjP+8xDNCcw0atXq7YTSZ39hSUmU
QxF4hewZLEH4d58sALcnX+a6WeOQ+tjUz4P0MTDVE+zuK2joDH9pTIGU/yoygibySkrwdDcolJz6
p0it69SINu5k1ilwk/Z7G7jU0VfXoyh5l4iNh91fyi57S+z/imUR7zT+OhQ48NeMkPQQMl2DUzl1
DJxcPInpTTja0XuJhUc3NrQKtJ1dglZDgdfIlDc75+ijxaKJ8LgTPm0ImD+mzBQ/ZHBPwPxyZ7lQ
y6CEqYhXPh4ZC2UYsAYlFCw2hUOZOHVBIBbegZBl1EGyYIkJSe5StiHS1w+4URE6o0Zw9msYlfG9
/4LyU3Tl8tX60ud4FzMxE+o+PEgMcdioDQNf/7CIr86jUrKv9QiTP5q/Z5kX3deRTJZ19MOJlnik
iG1CmFjXzCbJR26be5QdrDE1qsPzJJW7dymv7LScZVQ+lJVyr4PyePoMnPrZPuhjXoYoejqCQ82/
A6MOgN2puriMENx3HZLjH4S+HqIB2mzkxhBdUpUvXkRaI/7gS47z9pUqM/jPMOImS5WjoR6tqK1k
L40Jo4SxIqgc21Gy8hS7mrKYDtqLbsnv/IeE6rPwFTWvQ1nUlkHyES5PkDwU7zipONo8AN0139TG
yKjDl8JaQvR36twqSz4B+AF5Z+QqzVu9Tx0O4FDGrGPvVS4gNv3nfuPIC+U0VJOCXad2+fKQT2w3
IyoSSmcSokeTrrw4zCBwkOH62nEdV4WSRbsfsla/EpwYxJekjUkctkhDnYBu0n1KnTchx93rF1V5
LHnEGn9uB6yTOWTv/hlea9+PyEJD11UXDr0XBVFblkoEHbyhURLKy5j4uwNA2tpJAxa+2Raxu3t6
7XtwrC/W1zUMnmhZccKUrJCcxQgOJ51j65MhzYn8pIw5X6CcnrWmXqLy8NRm2oZNyVNhKqu/XNF9
FlQ6R/L/rbT4Zou7FyEBk3frhhSe/OMe7eEMuzM1Shw9QLKU/BEYjHJgozlG/ZIHkbAp7nhJJ8EY
PC1HzPn9ZNyN6ahxVJG59TloJkNZBK23oZVasTpgaWvswP267vKmrAaGGQuOWFBg85M+jLKE+6Q/
iQZlhEVu6xEhm/tXcMBiQ0B73Hc19r5sf8FNVOtuTPBCwYzXayTXeSNMkd9lBxQUkapoQ6kMkPCQ
tkv24R7YZAOs5Tu+TJsbsu9KE2UTu2MXpfCbUkVjMZULHbGTRFF1z0R0Qoyo/zBg4COSgnzXfiIV
lirjj7h/ze7HYpxvh6YgeezMl0WqSFAw6nSv+/hbyV1qd9sWU5TWYMw8UqknzTgdBrGwJmed6ALd
QIaZZJSn4Ph8/LdQ5vgPw7zqb9UBCqvFdi+r5bVbHi82Ao+B6+ar3yi0JoI1QaKqD0kF8ZG0TzJJ
gYZDMr0X2wn866IOVJukh11jKEDC7P4zaz/47XWmSthzPabBZkVZfotuMJlxTnnbMyphg5h7NsoX
rpONbpofw1x3kfM6Vkx/VG+JtVYaIr5G8vm/zhu4vD6nKbF2UxHdkPuHK/PD0Y7zzAY2qrYQdxTY
oFJpv28A2tQYJOxXA+hxDWv3oH2m4++JMpoFgy85tIcvEwQHWQDxj4jhdU8mOHwvy9rcnWDbwM3A
hFX1QgeGQP7gL/+h/2lg6Y+KWPkLs+LY4dS15EhbwOJOKiVlOJaB7aJKS0MHIVewoRdvvFp8wNbV
ts7j/wa+32ajnUlhPBT8cawwEUwHJ3VewbV3GPTk2UiDtMN6XtqEYv6hte7OZbigo5C3GjQnFu01
8W0gLpRjuUdTvmdtijnUJnujxEAQyd4pidkMIyEc3dSu8UEaj09bx8GghlSekPucnCE8MoOikSRu
eiqpxOuEyvxTf2p3nCJFyOeB7joxd2snjNCi+k+9+egdM8y8JLr6A0D//Vsh/7nBmbEdsizkv+9V
UePN+Quhy+qI8OTRCpK9L1REoXNuMwBs87svYcURilJ1aaV/opa4jk5ZF/qx4DPhcWbHraZhCdw0
F3VBf0KnZAuBdFSzrDnCDszv5w2uiNVDO+mLIWQe+joLS7epJ1802yRRE1/lRmRC4thBuOYpLLy/
1SAd5LrL7jOErg/Cpkf3726q0IU0iatoa5yKuul3MivQ0iTsdIbNl/BO2S5bBu0FwqhZwtHDTLNG
mgvYDEK7Uh76sdh94M2cM3PWoUKxXsy0M/OsIMsVUl0bw35hniZYg8sL/ACfuEHYAXK5T9Ykgxur
FnWHJil3oyOuqzO1kUV3f2hY7kQ6E4Bfhj25XORieK1yIHL2ZWxqttHjOTil9cZc4fYoKymn7QR5
MAoEyqfrsH8Xmwd7ibEPBowSsba+ZYvl2JbN48jICuhFwsK3+3rVPP+YFGxP5jvliruwMPD7s6hm
J5LuRy8CxIjB/ySkcCttF3BlUdyYJ7s0HwtogP27m3oal+mux+rU6KBxN9CvZFGH0IZzvzhpI8fU
C53Gtdte7cKW46SGF2+PzmNhlnPf8UDxsgoQXILvGRH0GRQfpxjM9q6JAekgzr9krAjMyaA7KtoR
jFNMEYrlHobCydaIM6fZJ1TNpyQo5+xaaUbtJmBhU5+pXdDoa0J5zENuXS+0BUd/BFIBAwfD5KaV
RVbg6Yd0wsjwcPKt6oP8y1cNgm431c6slHL2kjSxUiZ1fpBZX1FD29hR2Blw4Z6MC/IsJg+7W3hD
wnlPb0f+XXD6qlrxjGfcH2eaFu2DU+UsKpj68MWXyCOsbVM2fM77Pe/hJULHnygyG+GWfMX3abhO
8JW7jpyEUW3atndKl9jzQda9GYSHULTCjTXgEbCp64Qui8l8/019IYx68oGYxXJPf4EOFTaoBvFS
0OyaIrRbQbgmnLAHbcf3qFbbFEvfTNEraMUPMbGl7MB7KfWJJwV60Rohqcua//Ms61kCk0+V7qeI
atco+adGjzNIvmeoZzXFxWdLbB/XXugBxTdqlrt6LxMBCU6U9blnV867bvYxAnbaci6vlYZyVJn4
WiJ67c++5qOGF+SBX+VlXjPb8kSaJe8cYACWhhA5ZZCs2x+w+pebRRPJM/O7+2chDNBkYw/zh7+J
SQ+e38KrzHe1dl4/c8bvhe8Ho25ANVuPcBnBAOEHkrOA4hlkPV5C362cCroa/GNb9lVigz9lBWXm
vAvpTo0F68daDOgS+nH3xGBc87Tx7ZBRhbswYL38wYoLSnRvoNCej7+tvllzfiLR74car71hYuxx
gtzPC/geyCb/l6rkxRjflUYA0lQ0FAZrtOxlcdceVi5mbIieA6qJRYx57Fgf9olYG7XPgrCeFNfs
B5KmIpeS6jiRgr2pPGY4pbWxCaU1eAERdPxPs1BswHfevoS91vtBvKLjSOY/ZkAIagXpnBj0Qxtc
tCOUN8CbP6PG5hr2RA8AkjSZ3n53pbE0e/IZx8kJI3qeX/rhrp155LhttaopRQILOZoo4Ok8O9Rw
yZ1Bped89l6yow+wP3hbRdg9r87tl+87iCo8OB2uZXknZpFrPYFk3yS+RY4cQ9bFKHrJ2kF8zKX6
govkpKMy2g6HswhRMl5hcw97saKeFjpzpZ33B8i+YUFX6s0t1YvPBaayQYsmDT35kmzgVc28ZNhT
2pmeEF2EscDlIyIXqmOw4JOvltClRh1fDtx17E1nObkrwaGzUhGkuQYW8KAmv4ilz7WbtnYk0T2R
RabNrJn/EoBbg0FfvDtQjidFgthx8LxYQxF+PYqVDlrnNz2l23sMpx1L3N1HhRlEOw7b+k2G1AJ9
1HjL7SN6xlJuor/SQxRr/JPNXduFw7rHxGoNO862hw18aWe5I4T0r2Tg8E1jj+tvL4EOSr+Qy8s9
aVQjNaQuCszfih73kAcvsvFbUBRiqaX0moGT9xh2epi50APoDpfgxHFFsQYGsLHByBD8iDYOzr0V
tXj3zr7FJOCmpCxvZ5e5FHRKLRTWT7hiHR2Vr3tzPYUWhF7VkuLwrSw1qtXJ9LWFQk1nY00P7ucT
lt7CRupbc1cqqIdEEfI8jx7QJPWQrumf4OUYd05pGOpZaDR1vRGd5WleihFxwGvYcN9pXx6Rpr2R
zBgIL4437LFOl5bOg/EFLcyvYZywwkxh8FQW2Ipyh1b+PZoHPqAdQmd1MKR8/NO97oIiigmwUsrf
jGXkUBUCfUiGvbTFnjXJuW2mcWcmIRSFa7NKLtA6YWDsFjMdYQlAblDjoQTEIhDNQRXjFeB6Trtl
L/1IzEfcIF5dBPyNoUHM2KF/tCv3jSLZ5E/YuLV4Z3qWUfSCjRMGYsoKEXI/Mb6uXVgLTaAUDqAj
A+76sqexaDBGAFAzBLn+hlS8fZ/oZVxUmoSovTm+2v7wP59UAxwUGWUVVSOiPMDKOyWtZlowbJuj
vLnGkV7jaQlGvF6oDy58FCdD1yoBPKShOuVxJWPc4H48qbOJE4FcPpRMeJ4OWXLaaoJoFSXpTZPr
288eNxFAwiqwTgdeOnuXZVeCpZCSd/9iRHuiH6+aEVV6hASH0jlVWWTda0P81wMPWiRiyFtmhIWQ
gcWXcZxd10V56MGkbtVoDqotgGhcayMYjPt84twX0KI71ZifvAMC4TOekU4vp9sb8FVZPKxjfl1/
EnLnjA/I2iLHkzgFBcKssb4eMQgmGFu3QBKDCUSZVgVJtS2DkriWqDcArz4I32AkxMxhLiUk/YDf
1O3ZtdJ7+PN74apGCUksfHpDf+Cqw4qQmnzdtpKy/3rPt1/q7uyNWe6QlC+bWaLDTtMEoZbDYwVn
xYY+4W822U6ORtBr+0WMwbNRBkh3ScKwj0LmyRJOl8wSZY0gEVx1ii5/+Ht1ctW3+xz94v6WzNXf
9I98Qz00AfihwsszraEmlRWILUG+aO+UXaLzt1x4Ceuv+KMWfW0bxdI3o2X1OQH/WK6LCQHKkyfb
IFtG0kWaYVQ/BCScBGvKdNVkPhPKJVHHOBmhwDm0XlJq48mK+SJQT0jobBvje6h0q+fR2bG5NFXf
vCxiiIaDp/Xng89Tl8cbfMdz3RzVL9llOztigRWSrXKf/tCTnndDDdnntmknyCf1YBG4orfRH1cH
Hg+ySL8WuE3p+xJ1SDSpTTocXcZJUHc4WioyhhmFxYNBl1GjDyZf+drePPjDB6KaHr8YETyXMKg9
X+uKOfZInAYwGBZpoMGkWjoHK29VEOIMXjD54lq0kACcxK2Ti9I+3hMXFDE1SREMyRGnkzKoxKGm
flqPZKX7vYZlDXEZSwKDdcViHhUqBfSywEHA8RARVDRhkscQbgLSeYvWaBMa+pFmZDwA9DL2p3YM
QtaWmMvFUGN5ZIHnmRlnXyO5XlmDgYq0WtTGcXxEBVZBuAorzA2UgQgDgeJtsYPofwnxG0retxfk
7FTXx1aQocuWaXq6mGQdXOAy061LzJ0wtZvfEsWF9jBoqhS/4Mh2QKhb+OGoXHHsNaYmyWJqcWyK
rb1HDxf9i9/E2s9mMS/W0nDubzvjU7BnWX15qfunQ7ZRIAkryvzfLqJXSfpEbHkP0+eEM7p/3Ox4
jyqPK7HLa5sOD1E+scIDnLdhXksr50fgEY3oO3utkMNKzgKYmXnEv/U6rL2NxCusQhSJITP6lq2x
27TuzdLbdfYg9+FMcSj2a5aVvWZuC8AMHn/preQNq8At0ICwLZeLIqhZ2gFxiCcZlIvW0hgs8kp+
nCiitd1in0HWAURXR8wvJI6q1Iz7jkBMdQf3BCLZkSW7xHVjF7BoEKMH/83C5beh0FhmMgqwXeXS
2xT3EPOLKF8BhmogAYp6CbdEcJZlmBx/l6u8JzXiY8fd5RtT2ywdExL9CZRpD6LN26i3ZOX/Eqvu
l2G1FrExpQWoZqyQq3yqkPhlD6jzuLrApmR9yiccPFIDQv0u2lEJqFxCdL1gW/Vr6dOqRRpNytSO
zJ/JI+bggJhfzGRnieGQ/l6u839Fp8FuzUSWMJ1oxahUYyqMgDpQ+fdFmOxXxKHC9xUz3vo9RAMC
qydgxycW6AMatujPuvxBHpymVGnZJDRo+wAjY8Zk75w2FG2unfxttnaAn8+CKMezQjHjv0Ev/vhs
Rsyq+HoMjaUXyvyRqSGzFS2e+Bc0Wjr6qyeUX9AzY13xdgTJEE/TXoAQfgdIYRAftNfcWBvN5CpA
RPRLEbufQSHHSUzku5FbIGsU3Ze0UBi2duJrPycq8+NWwmLW+Gj4FrKdg49lthrJ/b75vTlUAzUD
y3gFbEZKR+7hxCjy0uJ55+ahEMAXr1e75TowIlwXa95x8qR7vJRqd/+ivKu6QOnAdTM+68U94AXw
2201DeyATyMBOiO6m5VpViRcpAXiAzLPDBwohC426Nsz6ppSi4Cj7XdZSyWLQvbj/EQ74acK5sYm
Rmg60nWfbRjT08jjVdrmt7rzFELpS5zIaom/v3amUqtzDw6MT8MXLtB22gVKqk2LZbdwbHYJLEU5
IcaJwhTwK9eGA+VCD0lgEBUl/udORqP6ASddLqG6C90Q/qnMOFWCOMMNTjD97jWdJalbS1t0QW1l
YGKsu1VoYFrmwhfUoMs2HulTfuSlW0jgcVlemxJFUq33NzEn0Pm/faoHrb6YPhjenwy21EwpDIQh
Ya8Hhpv6do1ekmVNsxfyVGsqsUGZ6laUlAckML/33kt+X2OlJzd/nd++rnbtePp8wHSbDE46NIgl
izJNrSue/+G4FJTLTeZTWQHKJA7vR0xyfDbHhVYWzXvsp+r3Q4LlUZAsotpVyin6EKHwyusliOo5
RK2Hux3r2IC4M0MJWMJ6kqCGoKBUZqpTP3fQT2CZvFf7bSISh8bbzzmidVRTli3OwCcWGo1BPd+I
sXQcQMvzTXBDeD22jzu76GCS5ilcr8X27VTksErO2TWdIa/T7BojfyB1UdN9reSxKwQt1RW/ge68
tHFVeZOaQzfQx71UmorZ8uJiAJ8QOFTMR+thuWQm8DLHqOOSvM1MRUBrg7LD9KdPlT94x+0H/PDX
9M/pfQ4aBt0L4Ouhqb2io2CpQOVRxDv8rmLZ05JaXBaXKbCKISt42v/mvqbJ/RxLOPlAx7dy8gfR
V6LdmLUg4Tb4+zDtb75gYmZGNsgi/Y7kg/vGgVccXTU+42HblOm+jMHhWbvoVDrxedYbdSb1ID1X
bqxuTA96QvRVSglQqtEILhjN838PKBWSwjXLHlRUctKeQAEAyWeccpzQzA5Zn0y95aImByenOL6n
fcV1fpWvb4f8qZhD8x4S2RBWZfDrwm5wnMwosoJAWoptfhJNjGeoaO7KB+Vau817pEBZ3kh+dM02
j+GNupR0u1izcVytim3kwLUSCQyEwBYcoKFEscZ8lbIUcZ3VPo45ql5zaju0WEqr6Qmd7GmYnGse
ps7ydibuuePquxZvR2h9q7I2eJYgHAH+3m7QS6CQDoeb41TEcpsMdyW6X2qRCBqGgoM/2g0oTl8y
OFACGY5YG4mg/Hi4FeGZf8HjHDWv+mZlQn16gVmh9pzYyn7nyM1DYLXFMR6CeDri0ATYIKZILGBn
+tfiY8viDEQVy5O6Z+dIiHs5DH2cXN1Uj+HOor63TgWZnKfGW6M/4qlk1cb7P3+vgSC1PT2SjaZU
nLljhyzkkxutInFGr4GL1ZgNrxhMXFNoCPdgWZ3hsYeBP17W4BwP2nSNUrJ0Gjp3Q85s+mQiw9mg
zqLBrWnAT1xZD+ZSZCFBg1z3Yo2IywMS4GmzLXzpwdhRJplT6DQ/QwIoCGmUbU304xoR4CnuAEAL
DSe9fW6PygGywNh6hOmPQhCCOnOHUAEebPtYpl7gA/6sk9GPyVKSnafY2tGLqwbLB3jd7hHFC1ju
NeYNJewWBJzn1Td5Q6LGYTEsrHHMlZQ7nQRSQPzS1FVrYKTgKbpjR/DR5ZqRzCmNRp0PIus/9ERk
C+wIQJaBk/21kqVKSye13rtO7HimVLl2swkJDRti5tlUNQKwry/wa8mmFMIfxM7+zWoABx8AFylH
Jz7qMtr+jv3Hh+1DbkNs8F7jvhbcMk1JkmAjCZqG+7u7aZEvRLmKD/DCuXhvPw3vDyWY5u9Inoog
H69v4lm0yDaim7/Mko1iBWZBZnN0ZLdfZsVl6TwY2HGdPhDFvRYT8HUXiFveSeydxAaKJUoYB3e8
On8q+9B7xoDfSI8Wj6QQUHqp9SQGnLXCkZ+m0DFdfyJoNrP9nUjKsQ7KUze+FREjcHswePjDf9m4
Gjys8Liy21Kk5fLAHChbo7w7LfkhfXb+uphzd7Fe7Dse0/e/EWJ1WUwc3I6U0YucDB1h6UgUqGpl
YvQEb+gZrLyzh6TbOxNJjWCo8nE6Tyo03jFz92u5EPPQP+m47iMBG1E3j9NxycxwTggp64Hmw/rl
PvQk5SHgqwCJDNii3SMn4a8gvj/MBRjrlEbuyAAgt3X0/L3qGsUFLTtT/vagxNEBKWtpiQ3WGkOP
fu42haqF2FqbcSOnXAO790TXBPea/YJTM+2xlMEJwkOrTY5M0hlwJk4pCo7r7zz1eIfTLQxajqH3
BgM8HtOuEfBtxJ4ihJ4fh5OQnnm4jbrFTRI/1G1Vvi/avs+NIJauMVje2CrfrTFuIYioefArJ4In
IeA3LiwBtVuzp5OXcRgPs5tr+6ox29OT2s5JyeXTE0lebNkkIXTGWWIETqZ22tspWfCPFL+3QfMN
Xhp2vR+rrUCan1SCX8LxaypwIXGCtE3EUJ2oiSvpRGVgtEYdGwyDyWMizEA/+X5GujqMj9JXCHfv
mlgNPnnIiT17jY8nMsl/dYQ78vvkYJeWZQbilhKI0019+rBDAKhNFDj4nwRk0LX6EUjxufTVymF7
yBe6tZzdAIk8rgjcKpG8f8lCiJ2KIWV3epHXHidlnvsf2PwH362ENQqM9o3AgxDZp7QLFT5W1Ier
NvMkeVklVFXDA4UjoIaOt2Le6r/JqE+65RRF6Le4n6h4OFOT5DuP/jbtYOVhjQ9ydc5tKQ0mL4WE
QthYFBYBJjazmr9MCAwATR39wSdwo+Ekkmd/v0rVl6pHsZV4PnaqCLz6Pm8jbG+zQQ62hb8a5k0c
51oKFgbMxuRjtP5OYoIPVlL924T+UsRp6xH1EvgYRnxMMqHilTPXNK3yLHH+w2QfrHp+vzNdJ7io
JtmA63gfuPLD74wpyQZ/+Y03yOsQLMoixSPciJ/iNPJEu3VRozAiWCvM+8asxkAQLte263+2yFS2
bMnjx1uzRoQMN6Dh8Gf/8BvX35Jc3SstfCEoB2ch78XjVa8ygpQvofdpuWHLGijqbsUJGsgOJ4Rs
BpkMgTGqP4wmeYZLx9hQ6qv+Mk7S2ojMJwY8ouudiqD6ezHaAXWfe2tdRg7rWoaibRb3UPk8vtaH
O8t0wZKdGW2p3wj+vY3ctmW5hJGWjtr56tZ/4tw147fS69g7hDk1kl0QZXyNCMCYsokOgLCZh69M
6AyCQpZsYECL1lBQYQWv8mM+tbhEDQRhpxg138Ht6PR+XnCY8E+IauZbctpI9aF1gY4ByoE5trV3
eIEcafoO5I/sEBu433DmlBg68Z8FGDLQBiHQX+iwUGiShX8tSfFc3ke66B8qRVoHw8kbbQFN6fsG
59LJf9SZT3+W/e7q/DiPf/0+IMXLHRfMrwYN8m6aTi4KTv0zmIdDQ9487BCiF/xYpBEGGUx6Zw/I
vuCZsNCwkUtAh3OKAn8gCgzn637JV3vwWUbecAROJRKPXqJPbLnUydSma2fd14c/0gs/XLd76Jww
VznQaCJyiR5n/VDlmuNk2kKZD5fWvkClQhgpqa2qpQSVT5DcKBeyTXxG3zmUtu6B6ofN0CdoBUFM
IsGiSCPY+U8E9mH3s0i4Np8ZLLvfn8w+joqYsR5BkLR/5vOqiqvsXRAXWy94bvClktcUyfOQICWu
qykqrldghEEkZjaiH92eoKWRDYp1ogH8+9ajW66EdoXeUiqUdfsS+JybiRumDZsKbI9yEmWWmBi7
DUEBHb0QKemQqVRbE5I7nR3ys+Lv7leiU0ZpNStcytdCMZbJ4KqPgc21xrFZrLBP9R7jkxKCgjZl
qDxd3tWkGYm3vdiELb/HC/hJ781kt/COo4AZxTRUSJv0izJLlyPOYITSOVgUQzT/duPV44a8DwzW
JZj0upObtX52sChe/rQmpg3cS/cRLxa3A8I/xeIrepUob60Uuv4l7Sv/JEAwoomAQiS5WrDPjB+V
8QzzOOwur/RxlobcnrRkZSvZytv+62G9d47+R//YBxaVcVIW0vl5Ora5HxCcZFV5npkc8DicjnQe
pb+fh5JB99YQ6hIw9XFPA70PWdYMBkLwRecRaiziZAq8kAW+tJmHrcCyrGtC+LXIKv30W7ej2aDm
vvQgFM/8bWt2oQL/9nXmz1zOBAbKptnKL+thnGF8xmTxjN0iEPfuGwLpCbKcVl2+bhFRLlb0DfEB
FmqP3MyfapRbibYyJkDQy29E8sreeA190ekzAVQM3YVztbiHM+n9zIhlAuSUo5zFetv6AO/SFLBv
AN26JKgABAuekGhyFeDqgVu/+43a3bcUD/o3M7tnwlLMdG44tEbDvMun6VkeqsTnGEgs7HPZu2gb
SY0rpYRF05i/7jbdC++Xoq7vnJHGDfBhkhhRK4zivMsKjzi8wcCvTy/O/dlaQzM2wffnutNjMOvd
tB29A2ZU2gtDPpl6VdcNxdfkEvmlLbFWF0Qz/ATfYH1u8dYXrVrNIZtjO3zMeYcmkfvdLpPzpVqJ
KosYtSyb7bSpQgxRzI42FVXeNTdXEz1CnkyU2/JbobMhHdind4JLNPpEWQf56TLbmFmJDtphzNRK
eEFvki9xn0FVD1id4X0ugX3IXO/aDeDRmkH0FLkZrtKWU4qMCN6M8MfgjfqULsITkuC+fKPNGzmP
aKAs30le+aTNsDCxq1XcXu8umdS/HisD4+QswzsPP4c1opkKpbQR3DMwkHqBDDTVohK+IP7yLp/T
XfAKVUjjOkz9h6EBlh1csJ9GnO6plYBNM/jFefq4Iwp9UgkzLIar0nR2u4CzobtQ379B07YVoqFg
YLFB/RhkjJ5NBB08N9x1e6+fLO2GbvLZpEEf1SSpy2eJUoL2JQfFC9+DESQJE5D4BXueB9UO+6jc
uWxgkPGxOi+RKuTvN/J96W12D6fgsx8+zYgcdDLgwSys/lOHuNdhzgt0E3pTgewaMA9Vmj1dLtwn
4xMUGyIGuZvnYCxY57dOa+X4k0871cEjTuEp3tEbg2kKcLjllQcv6Yv6cUWO8OzxW935i8/jwuOx
81NHYhUQkD/kVxtFk4y95UPGL48ko6Cc4CpZYVWk3R5VUGBGQMv312RYLakWkOXoQJwNZeJPg84U
DF8/E/jbxQY3QKdF3HQcfy6qdF87uyNLZA81pjyt6xBOIjIUO4yDyAguFiDCQYYGxE+yjiX/D+sW
L8G0gHUT6ywNy7/dDWQCj5yBx0qot5OegmwkPFtgAsYAzUOVOP7gIeOyuFMTd+B601uM/F5z1lxN
LsCt/wUlWcLiUi9pU59c5FItsqOuwDbnPnbByWFbgIRJIRqsumFpZ4INFcXbLULJqdj/kNlIBTXu
It4D3lt9F0aIwiMnagrsZgyA+LopdBl848Kmy82Wp1fK+YxfxkWwpeJ8LispkAioR9HejwoRkwCT
2r7QpMYJrLlNW9VRayxPHJJe6Ksym6M17XOU63aZr5ep5ywF6PEE15iwDu07HI8V0775YnX0FwLI
9O7RxLKwmbscsHn7Sp+SncG88UFzkLrfkZfPpgk3qO2Mxoo4FmgFOwvM5AuksM9i6/uw0mtkkNJS
NCPZxbpdaZgn+WovT6bH1nwGw21D7rqG2Q/aBojPvv0mE49Lqdeqp6lp0+yT0k0B6a8YN8Us1vRH
gDC0iCp0mS5FgbWfWWd+jYJWrcZPkCqXuzW2E63CKM+nbQm1C77HBHxznS8dhARXK8TXpXXz5MM4
/EXzSSUw70rWK/26L68yNDkVN+BqJ5nekO6wk2U4gNjZxo1vvqqu0MpSQCQyezUFZC7LmL65t3nO
uFlQw/YYbhxHF1aqSKVvmiIrXl/pFRgdCmgrAzQDa55IS8hxF2fkEiaFSICZZS5Ww9i/Axx/XM1y
HlcpETI8CS940u0OwARdt96osnMnEKmFhOY/8zAnS+v+mWn4+AwzUjaGqS6xvBJQRChTsbdP6e+Q
6l4gHckNx5UbslwddJ/925H0Gwy+gg5PtdPJWWA2Hgzum5TjjbvJbs5wKchDt7tNLGfuqdaLXAR3
NOX2C2KUpmOZz+miom4uOnmxFHwSXP03ZOGqSUZn6efaWuhZmJJ5aCWGVNRHUa9R4o6QjtdSTzbA
D7a+Ia6Qn8HxossfoZRgVprxLxs2Z3RO23ahsxmUAOWWfaV1n8Bc2xtnpzhMHgLdjE6VaYjBupqe
7nT7s8cHrYCu2EMLtMdJeR0rLJjzOX5aZF0rt3jVjBrKsdJGwrdA/vPtYHwGREYqkHsrIo7awVjP
r7odQP90Jkyeg6/tslcdWKjAFelsM0ND+4ayRk3s7Vkc5LlYxcT6BVeu9gZ0xHBDJuTgTEulSkAG
f6QjHYus//ui/kUIb4ap84ag5xAsSf79tHFTsbOCBWDoQPbgKwaFf9br9MKXSIIeHCNVMK+WaARi
uiDkxayuZC9Oen3f9il9IPJ5CtZay0NbcFjvjMIxoYDNNFkwrXO33watVHiVfAkBMxoGqFKQmBoA
zAKtR5TXUKgJTCtKLbzzR28CFuVpshf4R1rfvUECYWazk8Ey46/NqpdvWTRw6wCKiBfY1HBm/iGP
fmUktZraK17tZTTIX4AY59y2+RWY8L5O3J7Soo2h/A99fC8s0KbMMBY4Ctg/+FBYmX574BkGs2bg
kh5cB+68yhIcKCjcranu7whn0cqoAGv/K/8cyorJtfpskDHunWOvEfScCoaEqVAQDWREKaEGsgPT
Tm69/fVSaZV5L3MfDnox/8ZGg9UHmuz6t9FJU2batf3lhnbV8jd0rsPH0soAKClbuCRdTTiDrAib
D2c9Anl080Vr10l4ywqLd3EDq7Gg3iW5GFseiYRDzivp/1Ds63HoEE99a8ZwLPyW+Ic1wj2/2AGG
Hw+RBpqo7XGpZzv350CcsX44qS/LvICdtJnfQXGJTRrKm2xnCV6yno7wMnucjRbdzaRRljl1w4nL
UQE4Rn9EKIi8r9yUII7VqVwuI12cgwkl7J1Z6DqMqxfRlvzuwz8kNWGEBaT0bTLXEZ0vSO4mJ7qp
ZjrATAAO+3wNGsmakQYdiWAYdDDTqZxmBuhDS3hjiIVzHwDt1Kpmgnpyueq6oPFVb0LaQotFWkbk
FL7zOLe75vjwDIFJZW9lS9L/HU6lL3cJL2xz/N6XzLcayI3L6e2bNBDQSQRWHZ/e5mtHsPSAwfWw
MWIBEkyj7tv2RmbCNIH2Ow76zvyWmFRS7trUm/q2Q2BG4mteMu07EZaPYeNa2NkWWmH/aJkpNBX/
P/BAUY0mv5YP8NwCDsKFgYQzbIBlWLPY71OZorcaiBbKzA5rGL33S3n2Ig4l7IQMuKsIeK/E0uNx
fSi4Plj/8ZyDJNkhSTB+lF9A+YnatIL0zyJ62ik7c/vIFV96lYNIQzfw/OjA9j4Hw0wkYvFMM4mb
qJ7qmOQNGwBBqIikW1U+3ytWmy89RfKezoBy/s+jYfE5C5bQOBUif57GHFwOEgubM2+Ig1hDk3gx
t72cdtC7AFmgipPPJILWUy3Z0lVQtagRG+XA8p3l/Xt7K5RxOOGTzyP4OSPHA0QKkTKBtBFEmn/e
UPSAoWWLtQLwvFStKAGtGzbii5eYRzqKbLWnGRS/ryHWOkS9TDjwLbhQZllPcJjnUsgtmTZKSX0t
7bEnNMLRDwaqD9hr+FfkAZPCic53J/J/CjaJyp+T/LWX0TWqg2M6+wGLPLTQw4S9y9Xp6myeBEPp
uIseCwO0KmyRUSjCnwB/8dOECb4hfwToycnEXgH3NliGRM6SCR0/NYRsQioegiKLR7NmoYtQEMaZ
2tyIW4jYO6zn/H6Tuyz+aQ654HZ6jwRveUvb6ztoZ3gLHAkWGX+2oaXsNDmeZwe8/v8QKX17Ia83
9CbUXXaIHUuc8oNTjORu/fXgozHZlMvyPt9PetBBWEH0g4x7m0GwLc2rGjwKaJhckzJ7zG4+uqds
lkZ7cF7ImApkCZJ6eFcCht8W4WuIlTblADf7un1HAmJN19gnbhyAI00D1/P1Q0YydgmaFWA1V1QB
Bgd9Ns2dklQS1muNfJtlSxhfeFDmS3tb9WTu7wMe7iRvEyjXrzUtNVsNk98FuQwXmF8emCbMSSWw
TaGJhQLYP5k1r5iQxGPk7FVv9XZvTmWBAgeHdPmrZydQC+44YQzbKaDzCeT7UkYIxYoZjJkskOcs
MiEZx6PBmPqegwHBfLcOX6+/yJR5tzbfbb8zcPQ+86nPxmqf1z6nl7aakM+ozWG8DVfkNteaBGjE
NB3I8rFUKpOj5KVRSaqH0Upa1++cKAdLx5EM4yzqSrcqEKK9yV/KmhqQugrLNrcYp3doX8APzO3d
QdrGDrCSAfDF5PIWQYf+q/hbzXaYN4SvqonQ5dDMwiQG9lD0TfY/Q1oBt1tAGtPrkhwnWUIDp9dP
xdaJ7QeN0axP4hL2AmQn1TxaE4ZAMxmUBZ3gq+xgqnvkZWjt9I018tvyzPGXUMYdF6dzpKVJ29/d
rfiql1oA64nL48nbz4bF7i8f0R+DTzUavf+WCYL3xf9ZndflGiBzd+MOFLn5zvyRxouijqPh8pve
jklTq8eKnxiwRJazTo370ljdKGXgIVa7gMOgPBY6jS0PZcIPsvCsasIvw88gwY5cbiwEQhR+r8os
Kb7rPzcUCmDzoNcsRoFRzhQ91Loe2TcT05BKIGBECY6SmV36A/LjsT0fUACxeUW+9Ot8mUS4HJ9A
8Spv6QHtmk8eaBZu81UtnOxzNhy9tU2lT8XalSOdfZSfsRguo4NaoOnDFX/DnifCQNwKuSMB7Dxs
gpM6lYTe63V8wBItSfffr0s1gNS85MweleOMbg7ZCCCCPqZx4GD9Hr2XwzJ6096zHIvnWR+Nq6hx
KfICf+UDGm5E03KdlXNFX727/ibt4nwmymVollQpNLz5qgMqRlGkaNNkCESmctMNkapqT2dcpxz0
3ot2IH76mlZCIrqI/vE7fxEw0pGiLKi2FNCQz/taNxxfJp1Rp7jc2nNuvCCKvCjKV51UqR++l+nJ
r5iJUMWqGiv0TvZ0kiBsi4N3brphRefCrfeOMuGX1EffrOfXFKR/o41oYBbwSs0djn1+LDe0nYqU
DZ8Ny5aCvySs1cCBwq8OrLZHzwjo3iwJnQipsLXwbOKo/Z6evUXoU6EKWt73+guxt9JfB/eImQc/
WeliS7/A22F5smOLjtVpeL7l9+IpEv6PNxG7zFtC3fZ7T44J+vjjO5coZaWYb6bQW9gMKrKCOl0Q
NjVGv84GB74gSKGU1AJk9n4WIf0JEVarN8cOYU8EXOG3aym8bRfiG3KzkMDM7MS5ZpXM1iWjMrF0
SHlpNHLvnAoJyvNvkDv73hspRfyvserYjraMYLPrhXg5HdmTjXXAze+WwKIyckn8VPe4tx65DwX3
XWrEkZf73TZavdEy9ul8CtVodB15b5SXKFFIYpzjcuUrTWAdUTFKDMW4cso9Htp5ITq6Tx74VsSY
da2G+19SB1y9yISES9P2UbboCV/VL9kurFJVqpu2ltms7716vhXyv/uHvT0LO1SMpayV1UpGwVVL
aXLiVK7exkF30HYGcwlU7vQ7kNdgLQoT1c1qq4eJOXR2VRpbFY/53oU6TaZKH+Ev4LNl862Q2Ezj
Rajxqb/33tWQzSVwixG62o4r+2D/h/JKKst3k1bYWR/0dFX3VSiSd2DbZAi3jU67YxxcC8L5hVdr
QUjZ5IXh/NYj47sYGxJSJFlmViqHKEfHEPkdpCOPMmu/KpMcXNhSsQ4b7hVZo+C+udAlEzGvOxZy
XcX+b+6BRBIy2ckdMq8So3wdznpXeBxj49ebb1mr/tn8PCjsYER1n5zvJ/shelXLocJTVzv7A9X9
I56s4+F9hy0e7q4mAFzHVXPzVjj7NAZ52eR8lCJL79bP21h56ynLvFkdG0zud3xWTtI1RYS6QB9D
N0FfZjCvQRRwusmaoX8jb+ZHqukwjS/KhpC5X5tljNzAU6cQXB15jmwaj5VfGyU0LjanFk/STc+F
ZoYMiz2IF3f//Yy97Tld13cQGB1AUm8JaKWW7rrSMbJ4uyjxzuie57ICtwZqQgK1oQvbuc4VABPy
dtbEYxZYDv7I2jUPlPHYXXjvaE3JB8PRuIYMXkZex0QLl7RLm7v60zT2uCzYKiqorCm1RlFad/PH
GxsiudHj38YJM/podDJIysSbnoPpqSez92SHskfYNtv217D3+wajQrlx5/aceCdXCS2glOGOTEuh
jdO2hPvxFupxPiegUc14wwM0FmaDVfutYZ/BpWkYklj020/7E9T9scqe7jyWpMy3ys1RtuJqLEhS
pMzVmusZXmI5JFd1Kw9/e8nYrjCqq+roVg3vpKyDCpqJIErHkQOpMpExEsQQgj3sld9NqcagUB1h
RR1bGObh0qweWHJjaE35jRqRZRm2ZTrdJ7/zikxZpZ2IrSa+iz+4hVY/ptEwzkoCrRzwsQVufDEp
eIK6hcICQgnb9iRLAsiIeo3IWiM6kTA8rJFPRcijMMRbEXkapZ8t7kKeHsqTc4a5QoQh2Xzb3KHf
epcaTTXdM8IuNO5xkARN/zY4mAEmvg6OIIsJtpFBhLD5n40h4gNk+qBRdNsL47luN/ACN+/mxgXI
q2XQklLxUkVpD3aTHA7ZbLygZIe5boc1bKSB3g1qEOP96VoXOdE334vVKzxeZehMBDYCyr8vcJR3
GWQ4Mso0w35omucdG1N7DNoKFTuc3PP0xO58O8KgghkdFe/7hGtU6kfGflfum25nqokKj+4+yaBE
H38V0FFS6cbkDZDlvk46n7gRTDJ1gDvIPJ5FzTp6a/KsSbHzrulFsKwhXyqjmGBSIPqGvabMY8fH
WTVaLgkuBQ3tfuTGYOowqplhvYgXpWolFCW1TTKxyjn9DpIOg327CIGKqPVHVdljj/yf4rBso5AW
ZJS5wiU6j1dJm+X3ZhSqe9SfD8RQPCsfxpyMlRJPUAev2c3CaZL9nMr1H05P702XRbPBWStcQxgt
L5vhfojIykkNT+xUbgyLkAroO/QGIECjSApZr1eRslOJLJpP+yl5Wc9vl0Xv7r+qMt+GW0JMBs3j
lisKxFDGC5repoDBispwCcAeFPPKHg8ssl+a+2PZqy6HldmmffSMwCAIQqR5K4uDjAdg9uGji/zI
nu1IqLWDRd0xK4PQKi690hyIHKGZT4ZU17L1VI/Vknv3Vj0yzPYJ3Fv8HQv1Rambmg9+t/iq07bz
JxMn6xlYN6QYRJoQsWS5eMREZIBQFSWGM//+yC2rLchUWKVy8xielkW43J7Hl+g7ktpnf3mfNYJN
hzn7GEgIcn53p4+nsNkmy+2oWoR7I+kiJea5PfBybThVFdpBLVFHy8enMfjwt/ADrgi9b6Rh/RBU
K3C1fZhno7wCpKnin4Ir3N9uV96AcobfjrHuZ4quXl12rv0q7Lxk02HG4BMAKJxR4DtGqDZJQV8M
Qntr1zAiuSTJ9K/3nkL7sRp3lSTXhJKZdxeNuDRIDoVf/crkzJZM8blE3Hwkc2S45kqUzvSze+PM
dJWsBcMkAd92Zyygagb3UGO9PMjdK/FTobw3ZG7K+3tkRL+SmzpSAhK1QFhnVCfxgj7fu4R3yqbo
Dy1dxjUezGqBm9FXm82ij8EiWyn2sdZ+ce6XXmoWJ3ILBb6zHsCVSbi/V9yGGBgqYl+M5xoKjMWo
D6tFNOip+bJtPgKgRGzlhfPtPzaozm9WmaVeqnK3lZ7fYXbo4TmHlCkQ8eIK3cAUeprCdAFp/bM+
DKYm6wXGJ/TSRLNJRkXu5sfyCEF7IyK5pRVdiWGFZMp26dAJgzu9wt+NXFAhisRq643ggx8GOxfw
Dg2fBInTH3IlZpGrJ8niXU7KMsC0vrl5jq1H8oQuPv9dp7zUqMK1YCUb/FaR9EZDSmolrttXUXER
CZXUHL82XIwzooSXlc6R4kHAFUuBz1FEFWZ+1QKsKcUdyLuDOkFoQNTog2v3grf85JZCRpUBhwgZ
cm+PXCZdE5PhvSoyAgUYKMC3V7oDojce6pQsLTKcuWo5rCPiLTj5Xm0tcfEJ5q793LwhpDey7u+m
Kl8DlsLJ6DydHO+V9jNjVbujI1+Vgt90wn1L0XRHiuw9KvJuQRGscV6is/Yf3j0lthm2vL++ogYW
9j8/JDCkaSMbR21B1nF46unZS2nSX+8CLFrmTgHDXeYk+StK3uxV/elVZY44hq4fn0Viad5qgPW7
yc2W1j75XmLvsMq/wOP62DNsRzT3GHQlp15sdXXQe+jay5kZuMAGtqONw5xhTwoi8H6Sid1qBehS
mZDrgAoaFVsicwNlaMaNZKDv1msYuayYwmmJ2iunYWRijsK8pyT3Tb9mKHgyqUJ1J+NN/bh44pG9
zJwm8mXDCRts8TUG9TfZ8eXFmTPyWdS73uJVLX5QjT70+jMEHz5jx5AobdGIAA5PmwTCbXeBOU2P
mz0yGiIBZqi73Wu7M0W6jWu7ukpqPLTwVsWo6mropuv9nMn73lrHL/bsbvbJhyVYRp0BSC0Hd31z
82nB4DQGJ0rjjbZaWZLZCg7Fr1iOH50WbfGMTBjtQA++6aTN1Q6zZUiDJHB/f988Klz46KvTtBTR
M040t5yQatvgbFzkQZQI9LTGpoqRxvgv222IirKT/QEYz3Pu+xH4pRMcDSzLMHIzNsbwDwrTr12a
ogLMnFq7wQ/1qgzinJoA5G8PN60w/0cn5EVvWxctqarzNzQzDnmNcBSoPceSfwA0H7DM/hBvHGQF
jtHZNikqOxq4jaUqH9XedB2VFaAdCd3AzdPoB3FlQAYlI+6XysMKgJvXAiez+J/3THMne3KQYOs+
701piMe3KK732EAkeoANp9tGGwU7s5bX8n0L18GKzlzzml2JhgTWqhIDFfKmx2HZ6pOn+UKe/M4J
coVXKsIGCyy7PLfHxHbNNWVgcCxIjdvEjhsCPqtsCjdgmFuwInTdXG0djvZ81RVDxutW1mbUQvyp
ZFXDH6UNUgEQiTgXVvfL8p4jKAYlGCm4AjcmQYRL/H+5LAaG4JLxLwHc2nPiOh0S04T9OSeP5Q3j
ObkVzgauusjd81IQ0JDaZup4w9QLmHMw3Ug5fOZx8E6juqYEEWK1gStIKMVDCJaw2LjUT17QUHjZ
2xzXaHrpW529laslY7Qbn+u/RARgEU6Do+FlP1lj7UUSRbHLl7L5Wiu2vKSYW8mcnAMflrbrbmIp
D/kPN6RjAv5SBf1atdzBIQ6UU/ZhzqfgJcn5nMvAnKdNyBQVShcBggUKPYf6U+7Wmb69rM+0sb6J
1A/AS4P77unCQ+pBsyvDOX1b7Yd0cDaG5MuXsI+OmsD+wOPD8JaHDEsrCHrjlxTt8xm7b5oZapPu
Ks9c4mY1PXoz5BdXgCLoD/O8E9bA6bhtnB1L/yr6kSeHe4TgsvFH0nNekgyYnPoEofkbNRJzjqmt
SJWPbUqsDdCtIg92DMB1FNk4wsXz1zgnr56JlixCDa/4gJ9ChkCyxfJGb/NjOv7RljUEJ/uj3ZqM
2qJRnpWBSdo2Tg8+JBGcfFc5lT6bb/ai7kS7jbsMsMcWqy23HHbzwnKRhAQdoJYe3MZMP73KR/Tf
OfNmJ8QIEMUEB0P4BL08iom1HsyrDsrbv+3lSU2SUtElCWsdFo3HHhWrLjpMz4qzUZPljAlhIMY/
CjXGohun+WTE/RP+5ICv+WZYlXHX1ZWIFewMlyslWKgADTTlc1V2BxW2g2sEJSr2sptYjIQNOx5h
wZvz9xK4K8bSqXwFUzbJfVjt3E0O+BBM0W85YYykHQ5TZI/k1dpOmsH7kcnwvORcXPUMKUii31we
ZWmLMHmnEWMibe92yvYk6Q3lZmyxedfCWBC740pn34LaYLhBJSOdINFRoGJm3lyS8bDUIG83BfT7
h/3GcwVgXPbIIGPreFycqzfSBiRQIOfRBIwTKNfAb21tI+9uMZ8kMKc502j8VpjkllPLONV42k51
Eu29WEtwkC2zCcMsvuMnDxGUC+1xrJizLexh/O4VTQ5/itiXnoMzEK5PMdr3hOkISnMXjNHEc8B1
KJOx5HJwuT3Zxa/VfXCFHcdvnGEGGnrAnXz6YOj/zETZpd6bR5Dmn0Wt2fVKfjC6m78t32lbsz4r
Xl5tIfDYAjLQZux6xWB9dqZKF7wyFPmIaDvcMrSENVVfr9e9DeJe9s30WUNU+s9gMq7xRLZBEVqE
3Cns3syEgxwQvAnVC3SJa5Ruy4MOyMGclTwVWEMWgUwX/Z9Cvh/qEsfbiRa9YYJW9PemfwVXfGk1
ItqhbOPyR3KO1m9xCqM8gKhtWcskM5zoyPYriqbArDTJ9oJ72YtEcDZelzE5GKDewVih0g2tS4ej
hckIjLQUQnZkamJPJnhBjWN7cFWf3FodyUsIKd2d9VBYgOKI1P3TLrwNCVVGwKfcOHyTyxzo+9GZ
CkiaZR8as8GdQaYbqpMfAdbOcxgd4JYeJB/NJnoOpMx92hN+dTXE74RJybHMODoBrDFfOaCbWGcO
1eGvIcGArw2VV62X9LbfL1hNKNpJwZkNZVV8DJBZ9qJiuChGTKPIgs+/5/iWBjDorfl7ZBnRbUSw
Zmy7ZdRpZjFzEYVhE1NMycXSa+cr9rpiPGJAdTJixxc/Ojl6nur9sM1tjetAHDtGAvr/wYC8F5wD
OIP8TOeIKCg8tK6fmC1k4cuLspXsvEJ7+hF9p+6sre+QRGbIAudoj3N5x9df6cwYcoOOlBv1Fg92
IrC1kUStvkEOO5PhWIRgFLeNq/QrhHIGWaYoZcPKEeRsYuH3MTxiPnfdje1MqWtuBn3QI0RGY/kT
rrMMN71A9mPGW6kt7bcEu9JZWkNHXZNZ1yZ6CftUwtSnVQatjjXx1UUOAYBPfjO2WOXwpwBak3mZ
ox+Jp83j8T2ZKPWmxoUgxrrOUdQGtG1PVC0SnVkUCO3Aa2oCWuVaUm4OisazSomYODk+8lT9742+
y92MFUrntTj8L/r5GhilZUqE8xa5tamHvkz2elD/eVw0B+sxmZi4hGxr3UgfKceb/b/OT2fBRl9r
ITyk45MDm3ctVCbxH+MnDFMo9hGlsL52mFfrjWXYdpEG9u1Z5ay9McARZ91BHfs1Y+UtUqMHVDVg
ymNg99gzN+5um17lpk5hgo4oR0VyYNcDGVOmJ7IyaXRuEwMVnBTFMaA+9RppfKA/kQX7jRyfFTJy
iv78wfkEIIygomPgUfHzueHxIU6aHVfF3JT/3BXKVY0BSdGA3UijHa7RMGes3/tj2DqygsjPXn06
MahytseAmqxg7iVcCEF28UWLV30g3E9ld+/9NQARaefg0TYsgWeTHIP28pTGBnlrfRkIUUdJeMWf
FjprVwtKfVyHC5sTfpByxTfCWAOjgIICpffLO13LVDJnaBUXbxT8pveIZ4c/7XPvmd6j5r39tXxl
tMUdeIzuuAYhTtvyRlETy0dck6XB1UGLPmFzhecuDVPvY6lNjiITvdWgUQ1WH2A/xt5lYan9z71j
vRaebZKhwJo8QOPae68PZF73K9Jqn8NxQtsK1k3VrQVPLBwvidciefsGZ6W9A91yEMqZjUMRmzrz
qJ6pNokkkxV/2EaLVIX9R2qvuFoBo1txH1Zl7eOYcMxG6nZz0vysj2jSxVQREoZoB8j+9SpffR8H
kQNvRe/E4N9puV6Im6DygOLniUKfcNanzVnyLCslQruk9wnaHk9diUN2dSCI3TGFen0wNwhz6IMz
jjtu+6v1q5d64wRD1aBpflnNBQpByWFUPgi+Y0AC6DtKfX+5AFnFuRXVL6qjqrKkSKc3TdGd1wMp
c9zuPqdhYsQ29kIcLhjmml114esWuXFV9J0SkYATGZti9Z2XqpZ9ZfnWy3nKXTqqZ/drBg91EVt9
scnwHGmFbUlNPb4xlyOjtbsSfKW5nojp4fet8mgEqOfefrxn2YY5JiWKFY1fQLUZXvwVdszcOEyH
TPyClDVA+A3f96qT1HDavTSHTTkVFf8P4F1LWdKO/aXRfeG/+gYAVAq6xHPyVhfEPogGIlahvz2v
MI8l9H3oMa5YjYPWGaRuklhrN/KYalxHg+1kDdj2VQYTbzmZQadmyFhqFnyvWQCMGeM11Qwrsnqp
3e6awlV0PtE/olqHUhWK1YIfYGsW89R4/nnhIvbGMOY0WvWA4W5doEJLzX4ukZbyxez9S6oj2Iy5
BdwMX5TAjwfE2NflR/2Ll7LwU3SvXkSOUtcOVsEdIS+V9xqwrTzVLnNQn7eSr7zZLHoGMx4jwIk2
vTqF4aBVA45rzqm83ys5XedmN933z0eAjz2MpULZ+RacaNTgHqYcMYYDFvrL0Bl4ZiC8E7bjRJ/h
5IiDQlAl2FO/sM9zjDjk71UkCohTFJjMGNZ6S0CBTlaS05sRTXjBjE+VNo84FbpKgJO8ziNhouPe
MN2d6mAvJfIHjYlxe2cBgHSYV+/u9OE4BAao4Q6iYFLj31Ml1I9FzlOOjR8Bf+kL5NU1FdBkE7Wc
mlohurmqCO6fw9jdm31kHSdcHTZ5CPjjYNNdkPK0kYTPcfZ/tqXFCTA38rOU7c9zQUErluwPJIcD
Yeq8AATJlzSTuPWSHf99MCyLb8znjLE4yrKvWu/L4GaYMGDD6IAS2d3WubFMSBngLX2q2lC3K3hQ
bZZGilGM2iqiOFcx9SpeuU0LewjQbyfhZEY8FfYbN9ItCqFghDZUU583INYz9bOFIzhop6+BSKlG
cO2jvMZHNUi2Z5jZtxWZ0dyZ5KNJs0rWlB8/IWKIVpHxoL3xGdR4pztVhccFscZ/+vy3VnE2JSJk
7qf/R1NwJ6Xvu3I/3h3yM2gNbgBCqJWKWFEOo8PNDRPsIQR8qSunHT6GfFMbwGvnuEst0rPnriaY
RmmNg9juaL/La6FvCtf5DM/mhC6wFTLF4XcU565Wts91Mn/kbJwNlZ0Wj/WAGO4h0cUqJlqOEsJu
sW1af99dNj8I0tL2lerwADgVJkXu/KFCDelKVAudWmzzWC5aKyeGa/IunoVVKmYsv7m2Ph5OdM+6
vixCgLA8vOeNc4/P1k20kUczUCuDUtSL4UeDoWB8W1+2H+xw6bQtiBcf7l+8zrY/uRzGQuNsXAxX
E3oMp7oOU4sF2qT64pAE+EPVCxGh4EFh9LGKW7UdZgTY65FdpPt7le3LedsXy2vwch9KuRRAhsSx
QCORbMzyvXH6GT3Tg7EUEavi1/8bq+t2lmyq4lZfdCXSQemi+6diwB4RMktd9f4OLk6CSHwCj9RH
pYROYwe9lYHpOycb674ciKaJba+6OaKbCVo+uYs4HftAZMPTBJhSBCMefIQxO76Mt7krIYaBXzZw
jN7SVqXsATwjDsuDnCZlOWVAhXsRtDInvUa2jnotBcOedzQTQ2R+r6CwOzFtJuY4aUicjfTiXhsR
qRGE/sV9ZRpzBcuMLnc6gwv/gAVWACzpmgFf9llvBefwWgyjRCCLq7Kf+KuqxTVMzIe1QOCVhFnK
ZiEID+s9A0ktfJdnIAMye61I/znYEKrFmUz0NVJYmofG5J3b/bGkS1hFeSkDNphh3BnpO8791UDn
2QUvIeY6il5z4CNVHknpF/zxwyFw1ndNSIrD5EltWi/qX/C0GzMfua8PlYLnPwLEsIB8CzqfHQRh
mxFA96dYCdBLdOzmvS/j4DlyYXio8BHVjbiKvtf9ggsO+Uv0Lh0pD/K2CLNT3JfOsxEcQ0Gr2Zmi
o2b8sKy8Ld3S0Loli48xYlcIsSlJnVAkFjT0FsTxfAdzjY6eFvkRHubrRUYrSRzdo56eesx78Hoh
+blLoxZx7P9SM+zjEOTfH+PNxT0L5lshNX4zvaxgaEjzqua1hrPoQKhNpTBxQZ8Vf1FZi/+0ePDK
LdZ+3G9x/Zcs+FWxn6tlBAClaMw5vPQaJAgaIMiwvOP7gjHHQtOqcaJ21vJ4NoJyh3aLGzpH/tLx
636dRx2P4hIjoeV7+iBb1x6ysRNvLw/jBjxK2RMZ73mwzy++cvEViuBFHy5N4637l/DWZj2rPhmx
arjD1WDGJ3zfdpEuue1ybwFfOx1n+qkdSbT/SW3Bre8sVrvPxJykAQ4h3dGlnTszsARBHtrFVOwN
d6IpuBqFxJ/B+Q1XdrO3KJDpHnKgrs8vHlzYbGGTFLvjmIYwjfkx6xhwZVjxnn/NnpeS7Q5nGbJP
iYMZNQC4G8QKsIPUT1D8HK+5e1PUoWwMoyu6B2yWWp/F/fl8k3iKu5dpnQIHAlpQyvd2yuUTbasH
ink4PHx/0IAXkO86O2zPtOEpPK6thWr41HvDiZE535kgiasFgEd/X781piaXPPtUv2+//8XcnZ8T
3QO+JO0YalG2bZjH6nRzz9sykb2ppuodWHAL15ABwIQY7b0xabCn4XQJAOjjsoTanQBXpSR0BgKH
VNsBFdiFBq5/ZQcphsJE91plWYNNuzx1N2cNun863FUfK6PZrIF8LiI29xOdJFyo9dFPbO7GdkIB
B06O+1pclLgH8Yqi0BuXCrog/GmDFP2nPsJLsAlOAVGUQ8LyUzpMy+S3UWYDiLfngbbDyVTZFuiR
U1E8NRPTP6+q5dl3W45GbZsvbVYMyLIZn4W3wTgTGOGcLpZFvm2EO6l7mTMJ8QlNAbYDlDeNOYXB
BHsYxL0z6yyEIgQmpJTfQRrw6Hj/ezcEuj+THO3pA2BZjNzTQkzkY26SI8SRuazBC9UxBfJuFcOf
YB29mnzTekgnkZaZEKgxAoXSeD0//IHm/ot1kMpYDVXFS2LIaZbFU/p+/PW9BIhzsGvO6UuFy0g3
/9wmgXpH0og5kGb83OZWVqkhcGETDn9uKHA06uo3wyZmQ+krpr/0NrUWC03kugEPOzOeVkED0wAc
gX3kY8icltQwZBlqrvvUjwz6lTXKVqnoyKOh403QvmU1ncmDffs9aZEWjMuzgDWOhQf9qJA+I2Yb
fFnZ2ov1fkiD9xug3SiAiRwO+8fFCreEKOuOdWljBDZSFHSaGro881fA2/2l+QWTub/P4H38SEbP
IEKwYGJ/TqXonj4QwGM1uSJqDJDV5JsTBOKwsc6RsnMLK/e/iGhf+4sTaVpT4cR8E0ZVaZZYtM3b
lBy5/5kms4o5N9JDfDWFBp4+PbhdMfBS4zz4+ObF6ju6fWU8F8UyLfqVkNJfCuAofhs37DX+HRxG
Y0KJB1/tpy0NuR2zZosuQzgGmPt/PSFo4N/vkcw619bL0oXWAbeeHds83JoKQqsDGlkD6Eycq7pY
ga3cv2/H8esxPBbOC6a7D1Nn1xNS7XircGutcYqSU1dI6+qZmNyxiWHex8WLokVOzVGrA0czl0tg
Qf9mQPjIVyRuLISPjO41+xtgdbA9AFE3TEppGP6QThJRnB9GMHLdSXn/21AF6oCxWdumbe91RahE
8dbYpgisP076xfimMK4+ch3nWjSooIA5aO8RlXygV49+yqFJ4v20osuTWk41GCNF15aNwJoR+goQ
RK1TJ38OZzuAoo6vUt6HFYZ77QNAuDx+hN/lPezUtEgtqh0m+Y7iBegcjYUScL5tUHYdnm85tZBu
4M1szfATjlRtXu0mVTIYkyacpCVW7vzqCHBSKIbEy2QktqUFb/fOF6B8o0QKK99+ENeIQ7DSMNNU
eShNyXlvpcgmDcbZddWKtc1x6rmhjj6YM0/LYMUmfFKL//JKZyCQgwiyacOQ3O/iEOqxlBwuwbOl
xUoXnPOPXnczV+VxGCA5YRPeMhx4P1IPkED4+tIV3mMSietKAGc9Xr8/+sSBbj17dDA0SNLgu6T2
fv3iM0CHOMMRn6CjwGch0Do7UKciadYkGDqszQaYQCOiy085ScHriApv/5BeiIrkL0vlr4hIQymj
Gl56uxOq0TZI1F1f3bAwuTa3pn2JY+5WFLMVflFpVVUYrH6LS9PgBlT/2M5Y6L5Rq2C3qAaQs8m0
94rYGMOCp0cZNtiQ2Qd8zXqE7OS7EJSPTW8+wLW8hsfj2JFBJAj4zgrpduWZe7AfXHb9uchCWzWq
IXhNhqhzAnId44Ha5oC8rh5QmVNla5BBQEO28PqgNSea2WuavrAg/gusUZFE8Tq6N06E+xrZXqSp
Td9NCeHze5vJwfi01SG8cT2as2CQTD/EEdK7/lsXiSn9c5mArSvljpSzVDKOA/xMGPhANE1IKKyo
FbDPIZ6aWx9kS+lELSoL506GICa7eqZ2JNGkbq6AV/xMb9riD1PEQiiYs6fUQ+6FO8nDACs+jaHC
2EKnKwKj3sCNeL8QfWt6Go4FUiPWr9/oVr+gUlsTksfABt703I0O8qf27/a/ObJYnvdCY+sSXaCL
mnrkfLJ447EZvekA1cOzD2cPR0FL/HdUndyqTKBYqKJhpX1/6eDKZs7vV/+a3gC8fxjjTf3dXuUu
qgMIuPdthKby2lBkz4CsxaUGEFWKorpAi/Iik9G4aY0rOz0i3myifvobUXb8yWkvACtfmrfoH0gV
uhobuDEPWqDeIieeCi+6ScXZpHjDo/FraRCFV/xivJfy7b8yfDu50VxuXKiG3nb92hS2jMBuXz+M
zzgQWjcSvV5B0fGAkcptSicBmtGZSjjLbPYJZL1Lrap6UKAuqPCR7D7LIbVcGc7aX6MNnReFaBGp
WIrRHM0xPPQaDCkoYe7c4O9gLSSaxIwkZEUSkHTPE5wk72hTVun3zLbm9RyM7KuBS/PuPOD6NuVm
3wsDdKBMThxvh6Te02wmdlFvwsn7n+cNaUjVV/gjM6LXduZ5MjpezYy3o9hm96VRgTrEjtqQ+xNx
T+qZefkTJBbTXdvQ0ksozAIaKZKbI5lhTPNwLra/nk86hLV3iVy3iLfVpEeYCs7RTRmjN3x4fbw6
MX4hT1iu+3xCM2ZuCIgEzq57RLlcNyBb24hdfZ6T2Kc3VJnXYoBL/kqZ9ja32VJVHR8ymfWMTpLu
nnAplJG11rTMW/lzGibe1WmIJtIb02gwxDhBk6mYxjrPamjTBQuLsBifv/1U2HsUxY+AArFPN0lF
sw9JgYcCfLsHaF2tIQI2ZWfG259IyhvP0hHvwSX+30DmVpZqegjFZwSsWqC9yUliInJZIaNzT8GW
nlhy3E5JlnSHZ2qswvHI16ai6VR65SFuWG32XvzMWySQhsr4KiRcfSJehbTGLADdpiPX0ECYjqWT
2spM3gW5wduPz5fLbLt+2aJ77fx61QB3jJBa6Qa8Ct8+4FRiSdsRJymeoOc275ylzEa5L2d9M9Mu
BBvxOR5AjECQNGDi3PJ0FDRby594xNK/niH5mlH8Xfe1K0lTfS+3Nkp5dav4J12kAujnuJ07PTcf
uup5ItadM9dNfSv4qv/2beuWrfVE2G6tlolEPkbJNvbFd6MX+ykVVswCD6ovk00xn4E5usAfv0je
ZhogBHrCoeGdCQ1rL13B3rzhh3ZWH11j08wd67J+lDeyhJ5idFM/tQs8y4c28aEaXdV2iyrpX22p
RT92hHrhsEZ/yRFapcy8pt52hpN0aoTJi9QdXRmB/LzgEdVtnpCxFB4oG9oozFDbWhgkkI58TKhk
qOEtJRIL2MM7coMrtHoHLfB+bYVMtuHGwn0UFH8kYR/rUu6LPSWjgQYCjbDiBf8kQK2hjaCHOMmt
dmOYzrXjiQy7WFpwwHI0lPZjXDrgiAZiMXK7sgc0SelOo3xmewjMEU/2a6uhdjn0KqWm6gRAtNm1
qIMAAZJ0MUGQjP+izOoEOPzvZkGCEqSDxEgFRoOK4vCmqgBCLNGwPedve+OipImE62Etkua70d08
K2eHmXywoL4JgffFShoeY8NltEqR0TVwnKULMhuKCzFbtcbs2PvdCzPlEq56vJGwu4nLY9gkOCOt
3Kl0dIcHNlFqW8/USnnliM+JPPYxKsrTdc0IqkvXYJdFyEk98srFIT+hsn5PoNuIF0heMLkvbXDp
58wUKckj37jEwjDKO90fShSc+z/h4G2EJ/bWlGFJgPnPKGkOMlc3bk21BmVSMDBVn+9c6Ya+H31N
AdpUxzmFgZgVav3btVOioyayU9Zc5yZZr6tsZ6shyaYwD8H7w331rK5sDBBrMrLF1h8DodudC1iN
2y7zFVj6TTbE4q6h2Axk4ZaDmKsRL2+ZuAj4pRE5l9ZqWdHdyhJk9daS9brca+XKxAKln/vjRxgh
7O2sVNAA5kX64ZS3KWWjV8PJ+1ucw3g6mv3s6oW14VZL7lvKq4jBHnVsQZBfG6JBj+NhiL8/QiZB
gXPb3ofOOBek/Vv7xgmr2DLC8h4TGZcIZKc6gDBGPrhZxYWVv6A9snTyjZQzTnSKpxEjYOfQ8FmX
3Xd60MORAne7f2IF7PR6x4cgPEIRQYJxKPCyojjQD29CWHWFKPDIRFHwNVm2KeyfavrDSfGfxCSj
3bDovwMVsQZ5yV/X2NiUxTlS/R6HC/bkI8a3lY/a9wIS76mKcWal5sFaRS6t/zRpaHyjAIwiy2LB
M2CzF33ZAX7qy9rp+3T2f5qMsu2WkT7a1OBhLbXrc3kab/XSAnpGyd5g1YoRYLx62GeEV7YZSLp1
cUNZ9ITc7HasMvBspYTxqw4/sH+FGUoPVqZ60hCZexMjvPYBoAsY8kbwZyjwcUrnaVzXaa86xOeb
+M63c2KVTs0hcyInrPK9g5MKE7Xehb148RGqODztvxarYezMhwAHNL9Kjfrq/tsrsheUpztzkWMt
0XI+sSh97nv++7tS6YNNir1S3dYGjFxBot9FdPC3OJUgTgUbM7YM3yMRNvU+A1nYF6QS/Di0f2IH
WeWwYmWE0QKixM1ynoRg4TIm5gwGG+8/h8LzUmh4c07ECVkUg12ptoHsDEAx/1kEK7wiLWIMZUws
1wNL/vLGoK9GJOj6V6SNuN4kKYK16yAu0q2c4F7neJ2XytqPQc61Kag06YuZ6FOLUlK4i4z+a5SR
z7n9IMtISJ3xMk7BbFKcfxHcLRmCJYZLe8JcqfUyXrHFIJudxamDwCQvSn/POrUV6qZ5LYU7iCHa
0szcpu2smwU08CkZe5O7VSGH8UPx6xFMkynNw7qqL0OVH7h8C1DyHhXxctxnyOZmvIRtXtQ7Mixv
4KHhIsBSgiyEpHIVRyqVVX1UarOPZmYivzuqVVKEvtJcEKK9/h2oqWhn5gQa4LheSU9FnwtYUD9Z
+H/kOTtPDWFOCSovX6EN+FHTlLhirIu9FSREtv9/t4aRcCYO4Pk9GYJCcxiEfNiwuSCgpJZlNzci
mT+bQII9vGoc/zduUQBUlVUc/4X2x8gFyb1Qpweb8cqR4s+pym5u3DWPS+BDsp0RELC7xilcXPQG
GeeWRveOFBFRcChGGA2IJJ5Jfv1ItTH96HDg9m4dNL6Juh9OlMAthA2INjjgEhjFb9aU7Nfs0Up7
xP3uajeIM+335WmOxzluyPs5U4F4OX9cnpogqsmJ98tnz4cSCKHj2CIFsptoOE5rvnJR9SrSBCvc
DiaHacmEu8LwlWmu6wGwe0daxKGalvsgeb5KuXSwMJKnHZv1hJi0q/6+JzB6RY1Sc8hMxrtwr3jR
YpWkBTyXKMyweCOcgMH+ABtxPU/5ES5Qp02bE2Izbnrb/WbhtXnk05hQcRxpLtxXUTdTDDrSYl0L
GzYURjvRPR1X/aHm5e7Lk6G35uriDPVhKV4TdZHufC47MZRoOcPYgsdD7+Ep9/fiUeSHyWk5RL6B
QcVb45ScV5cHa7vP6YCrFghCLilH8mv2eJZt6PI7Yn98APmq8Mb6u2CbBZ5yD/tT/JsttCf6wcTU
jutFTPG1InInuEUy9glLs4qnbTXe8NIDG6VEPeXeAGd+7h1sOBNl/gQzjPN0pgcuBdK707+iL3DW
Q+2m2CHw40ca4B8rpS/4KC5oPEWG6YdDon+KUqW2uNtNrhP9qTucsdZzwn2xHcK10NxVV5lzNc+r
g/mbvwNdLHzYVDyr3oNDGAQMy4z8Mey4Q8ByYjnsXNMl3GBhw99cEAghmJN1gpa1e8ZSyRB4YTrM
ehBXHh01AbsY3nySvEiTPaD7j+B9ds9zQ8TfiZqFwiYPhl9cjNbfFU4ye2rNUhzaot75KKO5g0Fq
WgM08r0i4LXVYl01gsLAuKtoP7MvcZwJYoBN95Tl7a/nYKxPMcI1gB05urIHXpuNDHCrtp/SSGdd
hyl+nWFcS3xC5K9ynMpPfNM64udG34ACx08qP5/Z6XIxckIlgxiWS9bXScovy7u9o7HnCpbXnsxd
IEhKQAUVa2R6Xo/LAGqbSmfC3XcNSqw27H0chKpmz8Y4kdMMONyeVGp5oNcwt+M1a2JqwW+iFupz
zxXTD2Xw+yd/+oy5MGkVFuesY7cmhsgusLOky9n3GS8Tp7jopD/GEZSdk15fToxxOlpH9BiMKPik
w0zbiawPTY2FJ/lZ8qjjptDnuXPkYqZVrfPvXrkeXHoqLtEUj+thRxup+cExQXEzMT0eJ9wIJYjo
ywuUZxhyZwN0tOpkpVFkCWrZ0PC4GbwBK8uY2250YJ8ZXq+a8ahAn81BffVxS5BB5eMBC7GZ54Xd
qZAjcyuzpuUU8zjlSmGJs4BiEI0aHn+qc/5gHIgVlgY6FzQClP8IiaBWmb6ebAaw8acX1ffNhmFk
8/2PlUm5e1qdVpksLqu8EJo9EFVX61Au86afeiTHXjQIga5Jf6yU47TeIjtiepXnP+AgNhKV1jry
MLqaDIUIX5i5zJponAAF2Nl6X8FTHWC5hezvqLtI1pKw4Q00lX8F3oYqM6mX6OiH2J0M5WFldbs1
fKClX8Kpbm3Z3/fCEYCrBPuqcd/icp0GHcVire9nSQeCQ77TdhOUxSSuKxR6NuvAA2u5/0vwwIQJ
DuGM1OPUzoK5YR7ehA99ABPKujoERFXfzWrbatjbgar6t+yN/lxnUOqerN3m/wg0Zg9gccYhWBMI
VBvj2LdYo4s4xgPv3cbMdOfddYjSt1/tQ9TCzzVulXNc50m4jbujBrZIAwMy4mk0WRoGG+fi/V/R
8SrunzzYxhtLds3UdLaPxr7jzPDaxJlIHqHO4HoiZsQeI/tinhL5DTmEktGq7QYogEOheMBlseZk
sbaffDzemaY/f3q7wkIXr9UFOzNhEPNneoqt7KS6gCP7gx5pGpNUY0OM/rcRK2pBcQvfwUdjRZqG
/AtIRNu/hXMq+eB/DwQc8XJ7arYXb35ZfY4OUQlIkxxg0juNQQ+Us7W3qTfc9Wy/d75ToQjoFoKJ
SKtPAbea6WhNp2N7dERsE+vJUN93MPZYBfeCWPFMUhVfRAUa0VM/PxWozxdUzBqzvNEV9VAX49wp
Vyt3t7J9XcCdwRxF1NXY9JkHphyf5cishe/tnUHaVRrGrtHp3D7SG8hIrODH8PWNkA89u9cJ1n+1
YwcmuaeoaDf+SFE5u7aPuUtjp7sJx6yaIrBSsOJkAMlR1DxR/IpekGwuHivy8BxNtaM//OLtJ16N
j5Rb3rVrVCpPXsI37kSegOWtGI1UmKZIoZ7IZaX55f66VV2T/NzBiSqqLSBGHLDY7IS2NK5imVTW
C6qdXrkQy30+RaJX0Wdu+3fPpMnX8caqfoLDbRnuSiIBH4PqCu9blcndQ+i/AwYh1jwtSYF06GCb
Ock90qkqYX/TTmUbUdpHOWJ1RsrBEaSmZcBLu4t7ETMAS51tF560LTo7ZooEsuRHbo5lMHYfICHl
vgwP8hluK/lDUNhq+m468yfLa0KYieq++Rf1vS9qab19qJL1LpBb7z7QLnM9Bd+PYy5gheUqkK9H
beYVWiUzItTOdxnjqqR+xR6S7CnqEN6NeCt+NHvzpYha1v7gwuRPigqYBwKyqeGE/i1MpqPqCXDC
0CZrqWZ+zYBglALT+yZ5p2OrLOK+Dy4O5EZhwIVIS54YjoocucsEUKJR476EM/5J47Ad+260KciE
7QHC6AtPX3k2F3fyF7vbBqYnbn9XSlYy57B5g00A+W653NXyhArvNcPq7uh1Uc1UDLAR5jq0x4/D
o3XwEInT3Vw4AwKhVYF7PUnDJFMp8W9204ddhrLF0hpLzsMLIJ3yBPklkGlrbe91xi5IDCDEo5kM
eRe3lcvIp4udF5eiq/KzxUtVcpvXyRUTf61d8kP7jBuW9+luYSxGznIgyUl8g+ZUeUg0oU50mVNt
iBaxRs1kPrJFtS0zc7VryRU55iFDegR+cWOFwWA+sF/avzA6V24C+5fN8vnqTekC84JJcuJZg28h
ezUuX3+O/qUaIFP8T+Z4lBlbdHHZ3r+2q2s69ZUD20rlXBN3tsVoLO8hqFIkIQyTbKw3b7OY6SB+
4sKXOG3qhQldOlEtPRUD/HVejtlNl+nKbwgsza4Pu9JO4jHKoUchxxTkKZ+9YEcY9hO5AVXQJOhL
y7oSVhlnbWPJN1IbornaN9P51fvcwjTBL8XgNQoSF1XjMymJmOWTKyUHsrLzCPglxDraA5wqX3I8
RPIJlYN/4pPb/cW7GSi6IrjEYm6+/sh7bWj09Lc4APx/t2f8YRqs6WTkZaHgaErYgJATcNO0k3Nj
sF0hqJg6Etx/f2XIkVg0GTNo1/Dzp60blXM22+VIbif+A9G+pnh6kAMXkq3i/A4G+izBnxqe0rbF
0A1iVg+JYo5nDV6EeWnBHGSV/79W63s00zL8AJWOevlNNhT8M9Um1dm2CuTiAjSmbWck1Asm3aud
BOGfq8oI4N1wIsYBrBEuew1M0iQp1Lc6tsFGFk39GXQgp2VK/p0hOVhySAjWzZD5P2lFjRgWaoZn
QepYm3lJGrEWRJOQQLqMshYX1IFWvSN7SkD14vmSAPjQjxDDOoHyM5wgl5dtN/QPcPnS5oIbgWA9
AI94oKdeoa3A1vJVPQ6zm1VXcZOq18RX/b0pQkQxUH90ha9JAQMcLoGVXKX0HCESncBBQAnv5Bgw
Vv7WJVL+cBdQ+imp42GhvpQOp13f7W1nByQI+DUV7zEYhktPvNbPFouBTxYJ1MX3qDwX8aaN/Lek
qBywcaZa9pb8aZB3isdoMqN5nd+SMSRMqdNqxYafjdOTCOiTex0b/t92pcq6WuKr0r2kVZsFMxe2
GXWtQLTHnHQVSl18hEisIDRlmprF7uKwdHYmJP2E30KjpIGGw4KsrEFFXMf/5TkETvpvU5a1wOJZ
JpIm3no60mtnPvp64nfCHiAHlKq0sPwex25lfL5erRzx/sVzT8ihezLp5GyFXlgp7lMMYYgsc1U0
QyZk6A95I/9YHopCGzTtEBoNj/JnQQAS0LBiqykqvfRxLcxY1vgTGfQXKRh+gJiOh1mL/HmUau8c
u0gomr+VQwDGXDqG7QE4tu7TGAYqcOSRf5U57WIkS3pVQBnfTe/90IyNvycNO78ILW6qQhiwVVJe
i7y4a+gH1nNN0i+fVlXvXswxp2KXBiOOekii1J6o9eAxTM22WdkNWOfqCs9rl12Doc/qtlP0wS3U
BuKduJGoRqXlTE8rdTQ4yGzKiuLFvjQ5tT2AncQi96cBU6W/RrfLFH2n/7DC0drMQnCLxnitAfTd
nTFJ5DRN1XonTtSL7yJSKCm9gY8bTjiashxqzV57omI53w9ne3F8hdFxTnK4KV8fHdFH4C5+oLGw
Q1eq1YidPSMJgOP//zkWqqWZeYB9muM/fl9hCLszRuTHHi/tGksEYDhpR6MoT2kShddkdHfhiVtd
KdNdn1/RVIYaMpVELaojHsn0Uc71912BWWDyw7iqi2Yr57nCvMR8mQei9zi5RoaDWYagmN86TOnf
MPi9EyfWf6FbZTLrkA1uN2ALbrOtIA6YyadzGEDF5ZoyxXre18/goJnFyabAjzJjJoBroAMmUtr8
6zoWqJ761YT/MLeV5MYeZxzGCArOepvtPw/PamLjBH0joApGlkpcFfFk2OYG+S5o2FY+fjYmev/k
EbB/FPl2AF7QDZVDiBrqJO9IGtawfJTitJGX2Wvi3BJd1BQedKfWVLJr639CcYoR2nXXiJXzhJdA
Ww2peR+ZPAx2gMwVCFIA8JW/sptEbpzdqXDy9A3IGO9crPSn70SZVD0fQwUrOFCjNg0U+cBOF9iu
Nym3QzKOnBS/jIrlDsuUAhyVJKziGcOd2C8f7B7pIcS5RiRglrOfqS37UqhvRUu1li7thMdrw4YL
RsBSzlG2gIkLXEg/HtDIM5J9JAM8z+KsO4a5pPHS+XYiEwP324MR4orta61dZ4jjEAEZ2+BMMAAX
swBsDI8FW7p3bW8iM09MJsuPoC2EUb3bYdMOElljT6MjXK8ylVv71Uao4GIRSRtqsbpPSfd858O5
nRyfUep0yGWidS2PcLt29fQ7cxV0hOsJq94H+H9q/OVr3ncL0PdLh/+aQdDZI8ytYcCHNhB/tvJt
XXf4/PJ2jSptQszXWyUxR6k4Dx78mfTQjZqX3N7vwBUnL40+HNPqfNmL+7SlGlpZP6lANnJ6yXxV
eGtPiBhISNZFg7A+jlimEc0sP/kpNEbFwyL85o1RKiDB8ZoME9qcfwuWRiezNvk2rp9XpsBAPV+0
xV0GNy80ARERr4zK5BX08P96XCVlkhuoVZer4STuF2XgZW6s8ysHhPOW5MAkVONb2h345+AmQLd2
CxEI5NrwQlCjOI1AT/doHYhVXaSIofOa/Kcg1F0Aro1nzFkJP3d3ARk00AIQDsTf6C2U5ZHvyvhQ
O5XS5wuAGRgIwU5N10hxtFA5Yh3V79Q96z0lKIK9TDwk7g7aR1jYus9PzUgdMapyiXDfiZ11YKhC
eUJoH4e3rLV4Gq2W7AMPBP0LmDNguh8Wi37mnuQuKaYvSPUIih2amDxGsPVqq31461l3AJ47yfvq
kBfafYFsZOXgteDME0lVnbZUcazG1wxpkWpJa+HYce3NCdNsf7G8vXgnORr1puaNTR2SE8QhXTzd
5Yh90tNd788V8jT9Kyijx1ro9dYQyrYnXA/fDd0mgMiWPE97NiGuckRrvUKU/hyi4YKs+BP1lHXM
Rqo+4UCzgJHwHSsPAJoENXuNFgF+ii4FeB6vnymiwQDwMizNFc1LjnTmsOSQyhyfhPSplIyP20e4
DEns7hzCdWZckWYAPAWjgoLIbhnXUEqOmBPHt1+AwfAay6kak4Q3AUO2gh0w733RFGuwRpFfHk06
djlcUP9wFUBvGG+MDDTIKBIuKLo39eBHadVnC4/PoNqM5OpCdTaUC7D3QFUgA3LV7Top/OZqq3hV
pGXScms00VnHEfq4WdqpsZ+guuW4RYcMcwo9oDDnrdOcpXWpE7WkXbu3hnWh2RqGmCpITwaDbatI
k9rxc9pbomn0UJ5FfkRuk/ny0tEsmVMso+gMyb/pZnhVnOtiOKET1iwus9mVuzi7RUuHkc/l1mjB
8xLOUtP8GyZoDJBDFzdk9fRiz+9mv5NyiHQKKNhTX+bKaFB/tRpCYO5wjOkw37tBTPM2aTZmt4dc
qmu3bbNWq4uvCHKN/ER3Go9BuoEqsCuIGojNb6ELtWvo1vxjGRDqkKunLnLB/wClEUyeZldqwHzI
SxPOY5qQOaPDw9XQWtK5XYFJxIKcSpl8WAFKXJem3/ym4AhtAlrTZQfYXIMMyGA8WCkYkhfTr1dP
HJhgRpGqygyXghI04AOcuct+9/TZY3b03Wz0zlDzhxElm+VARJ6PbHkspLT9LY6/rWh+mcq6Hrhc
5lLmOGREmZDuHrK3RPoIMwa4RyzP9+SUPXrdLDAl9sLlPJDbsuH+camTLV7KaiWKZ9uagzWqqpbL
S1KTrouznh3thnsn4AfHv41WnZrTaSr96fDHTcnaX8C99k44eX3ueurlxHI6AdZmvUKSLa772pCi
KQRoGKfqNnpuHV3RQ27UUfYlR9+Yeehv4j6rswhLtn0KQjTVmJNsrsSu0pR3tTrI6ZyZZNORV52i
Sb6ODhRAgubgB5Ilp6/zZ4BVdVss5F64W3UKhd7esUMC5mprdU9ATeWz93+mLui7NBg9KiE570pk
ppaw0wxS5YCQtV5YMoeD8FSTHAvAfCL/pI3VIkeSKK/PaYBe3yNGTnGbH0GveYSYK7Qv9dF0QJgE
krp/EjPuwKaGMdDMZ2Z2izYLhAktVtodmfKpL1kEPuxZ4JMrt49bXtmynYHk65TSuhy7QWDx2YMS
vgm2wuPLw7NXTkHOGLHDwcy/Ok4Cz5eYrs1MefDC6lcPHwsDg/yHhtmz0rwue8w+hegIYymxt2hj
3EBavh477967aT7Ldpf35zgQOKoCv4mBo1Yx9qP1DFSBoCs1d6PSHoJL5xRLDfHfddvOd8I9UrTD
WvOl3CcbAmzT4zqpErFvdXmb8Ra780GyYz5SbW/u6QtG3Me+dDyUbyF0ehtWQT2PdbzOr7sSqCaV
L3e2h5NGuKsNIGvKoJz+l46quCng2O1NYQLKS3dcqY1ZsW2Vo7d2XLbbAcIfs6QZMPF0G2JYgbbU
Q5yMbkRsfEKfi5L7O3kw8UHX7S4ul77RF/wjZCXHBVIlhuB7AftfDLg+f7nhAGUwHm0VzenXmLf6
iHtog8EBQousdpeVBjY0uUhniIqVkqK/w53fPNXHgn38uM1IPGvLBbff4hvXtoITQjNnFwJkqn92
M6dRytr9MtirIHmVqp7G57W0S2QCj7c5REusnyvlVDJMXh9auEJjgsM4d/27exl8IWqHcJllMISU
QOF8V6q1oVXz7RorlhtDWfSqnCNUGzBZwGmVygq16L1cCj7rUpRJewvIGjfrGzrAgKUWi+EtjOKh
CMBuJcywrYLlRbP5/xiWe2a0n2Mhzwmcinmw/U4zlNHYNT8UfFaJyuapXRagwgvf+RqUlbi6PDfk
64iM0aF0AHULYLPh6/juDcgkK8d7rQyL3eAh/jAxa1vgoP91f1QUYwvYFrui7kQRclTfZ/JOBd8Q
ET6ktjUOyFwXZdPHaRystoS5isoNqtYnUNyS6brmyrSzDkrTDgQDFJZSFJdGNeK5ueMiujIPpE9o
VW3i3xbWxO/rIY3DwqycwQg07+J8gx2s2rFI8qNAc02IhSANrVUEwFruPJL3Srgga0CGPXL+wv/M
v55iKfbF2tiOLVHUZa7YlnKSJfqYkO//Wzzn8JJAYt5cQip70vJ0ZFTcIhj1LAh7XNwq7tNZm29P
iZ9D+1xh0OG6ZEjaoEasyG60IcAoBQHWo2KScxv4fqwG+A6a/+Nw9xkV3xmsJ10iE3gF8uXcYZE5
bH0xRzt+eqVwEJPPaw4+rWKIm3pkqSeEf3CApzV0cHTsr3pi2ztxl76IU+kSl1OiD5dOm/038p5T
vBlyaH3PLmU86cTOwYoUF5XRagq9FkAvVQDA0ZQ0yHkGqCXWmKMGpy6XT8q0Rklf3ktNHxBN3/sd
hWjlW/LeK8ZYb+QJeKVl9MQSZSNaLut0BGKaVpjxleaKZ2pWhfeNpvUTmLntp7Mj73QsHFo7iH76
moUpEn6lUvMgD44BsksKEq9CTP71a60AUSyzwvnlV9AwzgX9i/y+gU8cQG5GyykV7jWt9LSiubKY
lZ9shLvc2F1kLV+a4gOBi/mvaSEJU6ycNsIBxxC51795kZ2HoMihPlOdHPWSnwcZ0MCO8N6or4AQ
g7h+8QGze3FMeEGLZGOMICDYTU43jnTazeI819siOxIkb2hIXhJbNPg2w6fcRWFnuc/8DTnf11M2
9JkGG6JmZtEpvQBqgNk7oltUk/rC1ETrGymeABNYjRmJJnHVGVrvaniS2ALFOMzcZeVF0Ys38HoS
9urAywz9DDorVXi3r+X8CV35VOKcLuahMbrUl857JYv1HjDyJ7yY++BfEjWtQuEOTbehRrRooiwW
ycqyszajw8GFYRvWIt7HXt+qzCSG60wy7NliflK51koTWdCzdzsjMtaq+Q+s3LnLbgPquFIQ/Imr
HwhRMPsc+Q1P/537yCcZMfQEpZSGe7BkrQ/8Cbjs3uTw7pxAFsnr21NI2HK7b0V5bvwX8khT/wvh
/WVi1x6gHLl4BxwjmHyfRM90lraN03sF3O6SHbLG2WhSmgL33AgAqDTeZJQ2NKhFEyKOK5VzqFx5
18ox4vjhOeWWGItO5a+0lviWNDFqJBs1CHTVYog6T1RLMM4LvpkwOvDeDAGN8Nj5Tfn+RXfzOeNh
cj5fz2qnldgWYLE08FPI1i6edsbPMaiMjOWqTpe+xl6O34dHyPtdEQURqeq6vmW1o8tPTiz7LKVr
qXurfiJVYaK43HDyY59gk7+G9DQEo7NUuYNcvM/OWE7SJFkfkTQHWD277rY2Hyk+7s7GGQryQcYM
oyJeOVd7hrIebOxn6IIy9dm8fWJEvXnw2BhM0BPx67Fl7ple0kQrBoMF4jvv1+4slgw/aMSahhuN
LSFWkGobU3CrTwJGj3AnOyJnU4wus2odRQybhxf5giBW8pHIkLwymjnUJO/+mQ5SszI7+mur4kN3
GWgldJ+mT4ukvSRKE9BUl0RzCWHE7cgArKf+HdLePeekVxU5l6lL7yDVV73nZ8XaAaaPOGjkqBuz
Y3I7c9ExhwnDhwr1H/OiS5pzxPBNrMKkFbZtP/7YmDrxNwP+DbIz894dQ13vWh21SGIXktICKmWg
a++0GzmWvRJapzbbG3Tk6OlLI+iTGu53uq1v8NwuBASBi7apfvcRyevG0/husIaDLsBogaypUrQK
PAMkUnJ6aunhk91bGxPW26WLoGsFPPDWwUEwjxj6ZfDx1VjtZJ+VH2Wq5h4EzSDoVroS90jmDnxa
Se3xNn4uRjzhmQMlaCFgvu2sQpyJErzfa9vQlxd/1l5O3SSHm4Jn2Orcrup+G5BRFryCWqUEJ/0Y
y+EHOykiiByA+pz25vMAnPkUbjt7yYSF4ttNyhjwuICHwI5DJIbFGNnbJRcEB/Hk4FT2f/5HcNQP
HvShIcU6ERY+lO/afqVdTgfQ59XbEz1WKBeS/zciyympW6OIX0trdPRtW6jaCTUDSo0YdXuiD5h2
cN4i8DL5Oa8HE4S9XcGo3TuHFmIWaHWCII7w4IcJokVyET12cxi5qaBRlBTtcRhy65ZntfCiKz+E
ZwtNLjMSGaGqAzkbg6/qla3Tzh+90wsRPOuJY41auNxk3vKKgNoul6HgbFSAWrfwY+NGv+f1c7t3
94ynVCwxhvNFcYkdfXY43PA4W6ZMvq76WA0nuqfA7AE0x61D7j3G34niRILQ7ULOWaHRs6V/tCsj
HMGeXiot8kQby+w9DFD8c95J0CA8zM0Agf047D+DezW3QWbDLYyCGFzo4Ga3fHu2XKV3F5VTk3gK
ijJyf9W8QR86UYcRyWxsAfZSnhNwIbmrPySjflWWmyQFAsRgi0B9w+oljGLLH3PseC5Gs1iHsjdd
C6Pqk6fsLP6yB3C5Ncx7+Ke97csCDSlhTHOyHfm6lQ6xmATR7Rwv1EnfIGq9voRqKKryNQ4prMTr
Zb/hEpiVwgOCjEVlI2VRAfyiVvTbGYMo8FwWR9nJM2Ytb8jnKbVS4ryrtz+x9jieYPk5wd1Xrl1c
ubAMhnY/i8GNNacLMh9f6kvoGn42TNoRHirM9L16Mqm4JYBclYnD3Fy2Ie4D9MlF5LbNyhHNis3R
BNv7GOau/3hecTtF4juAY5g6u2nSWVcpBcEQ0fBZ8DBfN4jrE4GRG4rS4qPIE7fuNhkJTLIVCm/d
LOgsJihrh4t+/NdL4UTecSBWJXPZ3RhokIPrMN52RkXDwdNAV33wUhSmaDq4g32e/kovN7r65g1N
R8UoMJe4eQmsEjMC5Z71BOebTqXlWGnoD/S3hQS4O0xHqa9lNvritM0A85r4YspX4fG8KGqzRTlS
OaheMsiBHLwTw6fKoUvD41mYrExzbGjW0kV5k9wVyTZtTUY+WTmtt6EijHMgvw4pjhwDbpNmdmJj
5RMbiiIw9lpM57O1bXRHOn4/AlACssMX6CyjK+2TQM1wtl5nfkVWmGUuDz5wHTiTfNrEcqI1/MC8
uNPv03KVed2sRY+9Lh0t+kmuqED/b9WdANXmB3QeHgyjpNl6MhrT1PXGkYq57HkO+biTUKQ2lSwv
JjwRLstXzi9y2oGdpN0paUsxlZCl6HKfffAOd5CBXuWJGrEyLzcfGYqqrNzKUr6a3iqOTWFfSmhw
ignyRZ/uzKd+SOSVsgPcC+V9qjnvJVG/0bVpyEwbW64DfDR8AvCb4Q79vl/JusJ/wJJ7kcB0mioy
jO97L23O9BgTKFtX6aZSISlz6wjTcfmMIrGZoYUeWyoA2gzTG8pAbLi5+xDjD21S0TSfrck1mItA
0Q6Dwdjf2+lGyP/Z31S1+kgKeoQzGdQD8sdOJsDsO+XP4rg0N0V+A+Qp/pUktQB+8ZVGYuoCUqYp
3Ysvmf9nVsVudn3B5RvFhO53gCCZSyMgEAnJ5/BanUmoMiRiJKA1SqoO16dr5MLcW34mSqD7EV2P
hCrxB5xaQRts2L+mU+ziWInxYrzKH+35GQ2W4ob9+dQ44MToOG0bm2Qse5Y0ITGIYqOWz2fqS4XM
MmDB6xjoz9DMudrza/hqzfSPs8NUop+26NwDyrPeY74p3hsGA96RbDUT3q2u+7kO/29LR04+t4RP
PdcVYeP5PKBJbOtUUB/cSXaEQdRnMH8pFdfqyRPhpIxqQ1do1pfzFc4LEJZbulYm/kWCTRJKwmjE
o1p8KmoQTSFKFa4VEuXUZB1uRGEUYe79VBI5BtdJY2nQOdIdv3wN/B/pscbxnT57XUruUj4O/H5e
OFQjGIjMMOCZyet6my9Gjf4dBW6LmjO0wP6q7Y0T3D7tLtmEbHUev7VhBf3NZuz1epu7dQ48BJ0V
39x4v682ZGpFPZzPGDapeAOrqWd2dy+4n4QL2bz/v8Ju2uNCLKFCVcOX7n8SdFW+Qz7qUY5piWZY
/LVngHdsXnl7csMZgEBTGVsPrQtR2MueDFuWezB0iaSOgoWfIQgdqatYsYzLTx99hGp4lcCp+UA9
8Oqozr8EoOMv4/1VfzJlEmyYHgv3F23XIPPT5UY8RnoaVFsi2Ke8CojlRmpN4833+MgMNv9jmkKd
VdaeEX9ZfqhBxynXarDd69X0h33uh8EUbjD1QhuL01tEiy78mhUx0GBV7JjhUCr+TzY+dp/c0wDN
QZEetueTY2+fvehK8+gbf53CNvy+xSBmAMazCBBU79b2AYIDyOd0ItRZOq2Q8GHbfmdXoIGr/1LD
V4mYyLj9KMrr1+r0sNdiIvsU6kkzhgH3KZgoIL69vfB90eAJ4dQBO0arEHp9xUudJkQJpQU5JoW8
Qtv64Q/3mAMirmcP/KLGDaXpb2Hs2LtuQU6Yl3tuF5ttELnbGKqmKsXo2HLFmcb4q+DNhEary1iH
qhPhv2lsj2oHoNBDENr6KIp2B2+6BB5f9XdfweMDNMQlRT6rFb/RA7yQkPJ6REJc9v1kZoPkzeiA
a5tHgyr1txU5dEFwg6XY3xxHm0BBA4L0BP7Twx9UsviGtPhnARRtR54oLCKSe4gQ1FI2LSZhEsuO
3EA0qGCTHSjmgrSYL0JmRin2l9UEfJJljHIjw6wdZkGJZGx7w3vV/t4Q4MxwnnC3cYLI15C5x7Hk
E75MBfEVipt03+Lgvt6s54AzbS+UIwUIKuc0OTZwd/kHKfLNSlDYQgb1jqSRT9c2Xqrnnr3ImqRY
XitzJ9+9PKGRZyB2iLZz+bjvpVT76vXQhmfdzc93ObBGYoqUtT+9SSLDP7JB+0lwtv9kbyPEn+dq
gxSmZrr698vh2MggF4lv3hzHfr2Suq6M7RE0N5/+lF4GgchKy4S1fIzSh1xVDafYIqFldeeQbPr1
QfPRgpb58IE0SynGz5/+znR6VTjeoY3XmNIjluRldBUWtq22my/LGS6lapszgONwmnSIA5uo/Hi1
PTFA2XtlI2BprPCJ4VAbw7g2Vr6Fd7STvgWp/k6SGHPstNlO5NZyL5kMO4mzsT+xDlvZC4rs0WQN
UIcLgAPBYT5MX44AS/D8zuLD2ma3CGvPUPuPraXnXnbnZWZ+HTErXDeKzu/sE5ombD0idSea9xnh
JTT81QdamC9jhtTpBEUzpUA2qCxJaEI9eBLCtVE50K4T2udBkY66s1pui23IzkNf0P4XbhMu0f23
KEYoNdgxyuDt/iGqqVkjFUb+8fRAATr57167BzwTlKH0iYrCdohcRbgM9+nO13T8PGfHgljH/e34
ORZItrvf8wbNmrAwiDXfCMOLVJkGtEmPL1mQGpdhZbsu8urCEDuoTxJn/mZyMc+H+0KYSwwBSTVX
TGj5yx0t0TzVVuIjIo0RZRauvCjByxju5mnnzwPxVeQNXnB1QN98tsCqwpFEm9UEWVNMVZWJQrbT
Bd5XSWQ3VGQy14GFbTYz9/5UevryNUmwcN6rstHzrTL/qLQ7hsejtSDLDZgp+4p2MR3ydkAacsjn
GKC/R+U71fEpZ2rtVRr9VMsZm5c1wIdr43VzmXe+Lg8LXQORtPt2y4OIJV1+Svv03mBjjsttRDlI
9eZvHu55gef81eLCZ6zP45XRU4K2Ob5YZqFVlfqTespmphaeqhDrdq1sHpAlG8UwLJcgYhsQD1z9
TS53E406Ics8/7lHcc6kmRqSO8bGi6tIxQYawWAvUjTjWpWV8M9p6paUqVhNGwJ6qhyqOk5tnc2L
WYmWnNYRlwdorEt9eXrx4Jtmn66h0i7pU2JgR/iVtqQFjjIsQZrAXXEzGvCdGxTUbZBoddlo5NQ1
khr8D+DjfYOX1sNPZeEI5x4l8d9S/ZKifmJVWKY/hFn8X2pOrROjqzI8u0FIA85qNwpZfAwbtQ6n
OzW4iUj1RvV3oF44VRYNjg62h7sToaJonhQ90xgGnWpvdfGADi7peJhGp60YF/oMhMu5ZEHCykG1
kr3HmPtaRIJM67oY4bRfmxqiIiiB8HRTSu7eXZrC26kFNUe4OMQbx0QpzGpsix73O7jy6Xm/XqoI
/HaFLABBk5RzvXdWWoCktrlCCoy8bNr8f/aEHctyuZJhGFhxK1v+5FwvCt0ACV6Mto+tx0FY0wS+
/gpx1hzFL+Ysd8E0rYiq+rALWx1eNPGMcLf4GbBFSpzXyfwi3dQYpBDfwMJ/OQIWUr7Ej6IsrlNQ
NYEpez18eghSK6A8WM6uKyLQB81KuZ0429hm/XuW7/maacM8lX6h/lCHmMxS2lDBzpeC379k5qbY
bd84774hFs3UxIVTJKDkFncw96JDNT2WwF3FfNQv7Ohp1he/Md5zCgiSpdQtSTuvlDe6j5WmBBhr
iATcfve4fzdZL4fC8iGPNVpLZJhDYV87jmiYBfVuQxgWY94hksKbi/HSuAfvzMlGR0pdyxZY70cz
2vTnToSKDd4yK1UohmjAwDyxOR8wpFT3lrfwdE0nM1vJQz8CVwlMlv22SLfwX+i8HD9vRYAbJXWo
N6sNS0UQLZxBSkRH7LPf15c576eziPGq53g/O0U6GiQy4iS9IrZ6DpHGfO+EixOCBwCs+ttrJh2f
iea0u8ma6bOj50hOtD9o6En+QOqR4Fn8FHhSfxvw3mllai91kze72YM2DYgR052IKscNOmU+LtxN
+WfmMwbrLCCT6eLyIuuLGrKAzZWyahFDgcZnjxzoDFaqJHWVCSL3E1hTCXCY6MCwnZz84pigGbpE
d07zDeLkYxYE1YZfoQmAN1nYwLpTutwyxY2DsN7zOPxqAVwL9q+wZ1kuFhrDhed+xyNZPYmymTuO
3EuDJtpfoHc0dZxiZJ/ZGjZ14l/1z3ZZtnOw80S31LY3lJLLjDsYfk9yIG3lQLbVCD/tpQ6P7h5A
I7ID0n/zFFNjnOmtnVfftRXj4ttGFt0b7/XUg0HAgQNgtxdMRn8tdIARL4p0LIV9pBmNib0nG1F2
FkaQeawQr3ZNvew2YvZKqyell3y8xoXMBS5oFuyb7M190NZAaRd26vB9ULINTSz5+br+1C9QRbk9
lWd0rr3LdNZlb+jAAwq0c1HQpJRX3iYm1PpRo2bCrGCN0Y/zS+b4lXzYZnslwoIDOu3j6MH3/CKk
ytnjgEU2gW7Fjen8D0qRMtWV+1SGpIsbECCA6Mvo/i/BasNS4tjs32zs/BtyE28iS9h1H42fmeoW
Wo3bElPSjvqj1khc7gx+byfdb4KoLnSi37B8PJDJ2+iRjmYvJNaW9B8kjpakOc1/kWk4WKdVDW8L
CGGC8mLyFCtbU+RKCfBCBYPwJEsJ6BeFSVJCzx39xuRFPw/DZwG8S3c0hPev5GfL6uDPy6WkIs+3
OsDSwrDnh5hiSAzXmT4Qe/rsSBe5Ktwh+EFm4JRzkpx9BJtq0vz/t9iR/wElI3plHE1UmjdFvPHG
mdQjQfT3Qim2w1HwT8Yy2cC4u3MLU4Czhd8McNOrvP5WP+tm2naVz/RCgIdb6mfEMpvLfl753OH8
/EikHfpAx0mSb0DiHSFHRiYX/2R2zoowLaZpvNsfR+CzEgxkGBnsBaI3J3SGg5iy5YXZDk3BdzXb
UFnOUfxkhtfMP+tyASzJruCMomNOD6gnPlkmclw0Q+Q4oNSGVKQrmiK75kw6vmxTrAKJKTDNkfa1
1SdR/VkstFLpkbM7Y0yoPtPCmou/QlqK1ELEsCi6/huZ/mSzIf/6AesvDYTTyoMoTLuKeNKCuAop
Ml36JYmfnpyf4LLV3G7MUplvQ2FGGXgSkTrGOhOPN0k9nFsnM1hefY2olaf8IGfVO17p/NnI3QLD
znDe8mSIqYAJCDLwNEjkaPNBNXmBDEROIl/+SjVBPhiZX8sfxjY0puGOI3T/yakGs2EuGde6Y3kO
6tVpGXQudOZoPRpYX1Nj2/JDfc0SIRabd8+0gmhHVTcfg2pISpBb1eQ3bnY7BxASKLNsJ2fIIQ/g
DsY6Pq09fEbMqMkWLH2T6W6nnXj/DsihyZ03VpAG+d4ZCwvJs0VOlogzX1lAFBHPR11V6INBcGZc
1m4imj2J6JhckJPqvrxPd6mCbgbFzT477A0XKrjaFSIbqO7Zy41kurRA8hbQC5AvUfOBGc5zrTGM
75hLkkR5SY/LzKodeRTpPLfK9TSnrsXimURyHMluIBN1IMMgJlVZTeJjFVBS7zK1YTnGvtYMkC25
CyEACRdYO0RXXmg7EwWRuQ5S2Fq+ewInW4rSzTEgd+vLNLsR1fy6rX8hdbYsHEthNPbo618Je/BG
Yd3kQQ1bsY8xW+qjuZILZwZDsN1jyoenranhI7OOEOGV5Pp+6ePyBhh1Br8kulv+h+nFmhEdVjBN
Gu9aj6L7ut4BL2Gcm9OF+l8r64xxsfM/ArqPJxROVaXHPrsDgwmgF5OKLN14y4mByRT3T/P3tUKr
LYk2sLTjz7T22mZvUlB6gtILhk5sPhFz2R+oR9qjmM3J/RcZWxGZG/HfdVWTGbRUp/muFByl5pag
ymFpejd5+C4OgiPRxEQYsQjTI3G5F8PvbZV1P3XRhNYl+Kh7lWBXu0JMSf2N1v9nyGJT5hPXDPZb
/39ujTtQchXnvyOUYgAqCB677wPnvdqtJeYM3Hh2TZ0DtI/rlwwjBl5qqmWyrXgynoPWuy4L567h
67uRX21Fk9ETPfB9wcxd7hv6/ZTgFx8OWw1e8qvUEMUS5kDTLGlYBKybmB3eAw9KfhO3yDfQb3pF
LzYh3IGS9tiIyB/3mmBa2yw/Oe6mbuSLC1XwLfrAjTCLGz0yBfMH+Ia2IldGgv1OLnCT9A2sI6ol
zw8whpuETIGZe6Qqc8XUaMVG52KlWWbqnZknOda42ywuaczkTbPee1KL5JMw3FdK51EcJZmwSe6v
oVRU9W3CggX7pYL9wH/iVotZjt1l1WFZjkYRDThS3vVMyiIhHZKauS323TAuC1mGIYpotnHKEoQG
XFHFpocBU6pKTzttC1nqBHCBsQZcYQWxlGJmd+PSYU1BpkVX3KrHiOy+hROjOBXvnj3dMhMsiqCL
mkGMssYaS7zQDdqoxZuiJTaSSCSUEOcaTI7h+joXqzS6/xuqF4eKXpSytMZmXPTS8U+0L9549C7B
FAddK5JsP2Iu5MbmTy7XqwBmVFhTpBAtPOlUx8VdAfBqnc7Bfy/y+TrEsha+t2SCY+ipmX0N2MkL
CWram4o1HfzIugeU3vojt1wu/217cZcmXlbnV0P/BrDnHFHXNRNyAHeiTzcHp9GdU2BGk4bZz4eg
n4QKp5ywrns6lOmdVItQ0ezMnAQkC+P32GRxdoktFvSwgB3DAEcs7QG3W8CTh9ysVBDAorBYFO8s
97MUpdsaNfWM5R9HJYE4ekqKMU1z75TI250bTxT5lj6eLPeDWqwDssD+r1JVUW/jniazJtpbtLt8
juiMq12msOfz2yYsBtr4DuathGrnIZ4FKKgjAz480re2+jh7/zuuR46hDf6LxZzM6TNFeuLnDYnA
GlNSeihGyJy4u91WgqBxbENrQocXtedeYtaguRnMUU1VmIRSXU4fXgPH+JQx3flME1i8tFNV4HiU
fNByi6Z4JMSp8gdjjfXhH3PCx824pOow7ueEPsEzpBYlAwZTzoQxKWTROLEx81aWlavzagPBNzix
upI94wQYo9Pg+P8iyeWBOIpFZXEz5+8XcpTVgImlqU4aSnt/JBYbStetdJL0sbTar2d5lC4mNazm
LQZv2yBzVtffxHaCvXv40ZQmk1XKbBwmhDUGpdnHzTK76yQEP6DE4IFjaRq/vkfJWVVtqS3WXOkg
JdaPSVjlBtDBwQqtFCxRAGZpPtWPWRUmlMlhTCjmmDTgYMBOEkZyuhsjUe6vJNbewAUk7V8+3jz/
JLtr9zj6ZTOG1qNyGm4hGhu6qdu7oX74mMJTp9UWTtLd6rLMnIvC4ZS77HQG3v1TCztdy+jZP2Al
wvW6P+L84YbBNIOUuqB4U+6QeddobeJLmfq+ZK6n2XtqISQX1PrJQ9U+E5K1vgBJUDY4V0WogJjJ
LFTSyDGbbGYk+qx5iCNTtyurt9By1LlSuvwYy+eox9bSJpy04ovni4fTRhxzl0hCANa1uIpsn2Sw
RLfhoryT5i1/F7ZBRSHZL9XOvcZXxhZpgfBs6pZHZHW0dPint1W3sZmyAvYXRk6eFQ07UlafPOAc
zTGD7K7Bf5au3xuZnMh8gN3pbY+IdTexTLAgz7ZPRGAr2+PFUFqn2hOxaFPNh8139JwCYqzvvoZw
QAw90g86JvheH/NmYaiRxG/Ey+mLXdyXoL+e3g4fhkOtaFxWHRYMNTnS5i4LQqHfR3CxptGQobEO
Jn3ewoLqqBBss9+MNi6vmgbkxZnVlyOtOkPhaiEX9EsFOweKc3w+1eKVqwIQmbvTtabQpnFrWMBC
mWNE5Wph11Pl+5T2BJgjgcbwJXyToBt9cq1AJ5LtyDJyB/cePV3+jClDK5DRMmLsv16t0nx0KD4r
NRwfmQEEw3WSif3VeLl+oxS+oONYr7ugP4KNQGieq4d40XnRtwmhlUfYePcfJm2GmLYfFNUupWk0
/Axl00GyUb9alM0xmvItPuXOuQ3fuGvPXCx3jdZUfkwzUYeW3oFP0y0TJseW+8nAksRaTN+B34Cy
+pNaoSjvwFGOAZsa1hlaTt3BPky5t4iG6tbuhM7RUTLrXwUxJjxBVnEholBa+++IaLh6PQbjYu7o
uPpea7X0m3dG9INbiryJMHNmnhYXMSv45jVaWnYHlCeq9HuoH3z8Psy8OTjPeRIRHTL/MXmrQ0zO
9b8U72cT8TrjrudTeM6V/2RXRPmBhZItJpy08uBmg4qkRj+c2Z5vJE3+MSBlWPxYKVW86RjooYkn
ZYZdkxUUxmVov0m+pNOPoXiAteZrIiT4NYtFFroh8f3JVZEKgQypE7GMeIN5tozkarCEF9ZVuxIn
2WysiVoSUnm1lUtLgnEZha/AgCgl1dcRUDPgnIRKodLz2b6P1OTVNSrKoZPTGI5TL7Cf9X3aZTJO
nE4muAs6o8PC2/LCWr4pNMzJbx1ZqKkFx3ndNMKCmOt+qIqtc43eMld7R2t8VqQ2COLTKB+/6PXi
+AUxfRs7vG3nBZ14BQxVNNwedJojnetv+piudoXU7gDLvFPhj36aQMmD0S5O64KWF8YxkgQ/Rpbf
IjH1vvQxh9r7Tyfwi5dl/hGRCPe33+1BrKx/9o5101QKFbwLVPvzVeOD4znPNeS+qsQgC9msbl02
uPcx82x6rV8PPsLtpuWWn6osRamQk+21nyKF8EB6P3u4S0bDTNhqg0S4/gMxUHDdc9Yplypi8wc0
6lbHOFTul2VAm0xW6ieKib1z/1Xo5Oy3JR/ni/YsG9gXXiLQ3EHyYmQrqQuRRTDnvuaN4BMV6lWp
uGr60vmUfMLGLNY4eMwAbuzPkkY6g0l6wh078zNX9L0bF4BNhSrl8QP4xYTvVQ8coVaxP4hhk5To
UvTW0Dky9nizB8DDkGYcBBXS0eT4q1VbwLw/2Hne7B5H6zZRqOsJXUt20vCSSUHdS0Il9/mrGk+K
gjqMq3FXpuJCqJNZt75/OPpSg/ELUPOyaz39jJaq1gA/lPf1WJORCSptkoRF3vrgLDnaW6LwZ5S5
IbYd+KbBVC5AWN4JSYIPJGzbB13vUv+wqsUd8XXN0j6cwF6RWvnwdZ32gqbqo7kCo7tWQCwM3LXE
E5cT/0G55r+Y9wxBTePq06d5g815yv/ekYNpn7ctOq4+qrVi1B2PtfN++/fqiOcSh8JP/BN2EklK
23Z7eXOa66hOmZxBvXNYyQ3yFvI2HFLz+P5sb0b/aHN+7lZgPkfw/822EbrMiY3xfB7DfV6qspLQ
Nl0+PpmzCdJfgotgfaStZuMbrmhl1VGhoVkudOI2hQKut2NpY2veqfX2B/2NYeTu0KKc2jkiCIEz
Y61H6EYgp1js7PIkWQnq2iE2J13nhO5P5DC1arYODxEjoKrWBWyjleeN3k91jhkPovYMQAHO4/+g
lYF2MU8OCoRTMPSYlu8/e/HDIxDwoeWw0kVWZnePrkFW8Dk/A4PM7JcVLAk4w4jawAB+TKeOgPzP
HXgukYNk/wnr0+ghsH1SuBovGZP8wDkZcAY8A4AZuDVRx1OngSUx0zkRAL2/XmxbhgmhlPi9+sWr
2lhzNqOEYXy9j5H0IyHJQ/cqsvz+gIL+q0x+2SHpRMpsT/MsN1rlxHwNErrIJLu/YS192VmibeBb
mJf1WbH+8V/MXAkxwexzDsb4eJGJ7gPiNB+fguMhWOqNwUzUoTA9H6+B2GBlRJ1Ofzxc/MUYJzmp
US1UQ3zAQNmH+aa3S+ebn4VybMeNSSbf0WJo/fIP6Wxcv4LhvW8nmqtwkzspItDB4LYozLtNlj7m
WQ0ICco1zBx9s+ESakpC3GUthg7EP5z+LzAfjs+3r9ldt86bm1QB/etCMW+6I14dbq4XQlugOfi8
NeX93J5AgXqQ9bRdkP9hhkWEL/ZvJZUkdT6blKWm2GzZKFrIaEA4Os5cH+c721eRy0hjwtWJurLS
P8muJWQEkdKC8Wh0KJlmqs3cuo5VwGRrKBGcOnUotdF85zPKFCcQEPtYcn41ZWO5tEgAmnunPA09
rJsYELvurqqFZ8K0XJeU3vMzCpa9shSYb2gPQOHeeenTMSds5+iawM4pbAfic9YfnHBAwJcND+FL
3Y+/jsq0RMot0cs+Kc/QAv8y/3bktjs7ixLsq9+Gp8lIKpP/q6g3pqIwbDEmWWUGQT79ZnBBvwFl
jT/g6mMVh/8OwzzvlUuwXW4sUAWn/uKwsrk+u94CY1GH8YJYpty0tWDGAusKpCI3WEIdMF/8htop
bYypAPMG8ojmWQCAUDxaQSfjPh64UBp351OSsKnPpYaA6LrMdJ5V3HQUW0C6ajITtAu97eWrqAeL
/ALQlonVgzHmjbJdhEAhCQRRjOj0AefXsP0qt0KO1xtokigwHrAXp689+NV94hMio9AhJFJR3x9U
2QoEH/7Z0ZOkHMHjY+a19H9oCtVbL5eHQCUEckGvyT/TndksoA5cZmwDNhf7jc21WWzinPgBJyaK
8fjT4U8iDCJcYjVrZMg+ZLjImYM3vhhPag9LhbqyZTJklVLNxacb3gXt4joNu04sE66gGyj4YVb0
1oPTJr+yJ5ccQJpwDFqyy1gVJA+0JgN6N1CqNLR3Vqodo2WQl0wLexBMEWRrRgeIxVReR6jzOVth
7hsTc9KFdWJdCAJLTmfVcIuWbxrPZ/OHReQXj4te+AOQ7uLkdcJESgQubTmXxBL2gXv+raSqEU6D
HDNBcp6dNF+pFk8LVqJC5VzIHPeiCrp+SQUreMLmeTZuTlj5TCh5fmrwsgpJEFMUsbBWI8RRJZVt
/a3wSneo5sQYU4MknppYDnXWhsDnpGhII7rWY+Ysx446FICDQRxQkvfrOktFbyOXt+J/sJhoa6qw
LC7YoSnulsr0efR6iGchPLXmtJk+/4IY7v0UoWOt0QGh3oQu1qQK9n0FM+3+oXzC0aZ44w6HqZ/N
KqSt0ekVUfjZ9TYwazU5Th39KqI+RBErzxO0vo+oroZit9GbmCrXE0q0VUIJ71VN9zOnneOfcdzO
SFYx70TpG02fXsXHm9CxPs5SxY79YvWMun29MS5zcS5zuiobmae/h2M1wmyjRfiQ7FQ4fluxZwwL
tl81+iuiWcJiZhceeAHVbPb3raOFgTX6kkxdjgMk4GVBD7JhzkL8UHPrfx9o6DdIwR1U2C0hvWvd
yQ8tBU0uP77d2IRX6fjdFNsjE4Wct9XRL5w1Sxk8CXHGh0Y8wxBy2wrl4maskPwA+hCHWjbhIcrJ
rs5NWHlUUeVIGfdv14lRFIdLd03E+iI1hS7HvwaJgCJLve1XfBdf1j2XjPzyrroATiywoXlqYFlE
Oa2Or7MfVb462x0g4o+hALAGSo4NzLE9NZP6H5n0w3pWEOJSW0lM28tIynStovT5Ju5HylMr6FZV
QFZi9zPFsaHuvbxeTUasrH2FN8O4VVduJc6HM5k5JqrlZFOnj7SmcTEM3j1kyKv6U95az6cWH+BD
2hFPkqbXkEKjqVUQHTF74xNNrLOOcqzIZTCMCnlCfFgRowSyphxRlnZrMN/knJv8OsV+6EU2/UGP
UEkv+ASK9+KDj5ZFqBYqZ8uDTXWAhUHLKtJLUi8yflTUXR3Z4oydw0IZdezk9kIuBu0O9BLJi/OV
2k07cpNcUNCdTmghCAuiSmk4ddbr4pmZCHptl+icMa/Y8gh0adS7MpnnJK1A+xsTyKTx/+xxYvtD
dCoYcNc7Be5BuYbmyQg65BKhzwHBMrv+L//gBd8nEfR3aJ9rg6zhrWJp770nKlGOsoDxTHTZtIkd
Jf7xt5Xli4Czc/PJayZ5SmE7ZJ5+2QtHlERwd7kqXp0O3ksiVz2rk0nxijamphN6YWhEdHujNXzW
B7HUcDucFe8c2OqVV13MHoiaYLhy5AQkmQXUdogEFDVQZZ829lou8uxIbpKNSPmetJ733ih1esQw
9OHrC1+KkaZG8zxcoPshFgfxhzLoan+3oUxyKQMvedWKOEALzh/1Ndd9l7E4d9DZQ85goCcGbblW
nbE65KIz71zRl1x3ILZLGTXzNn/9i47+mQyH7Gj1rfC5e27ttf7r0F5GosHnADdIcx1+Si6EHaA7
3VOwaVir5PAcFMScAtz7WdktSdxqT2QGaaYEn6nNbSGoj9ff2x0eWuv760usKQo4dfhSIHpUgyBw
+0K0h3UpQiZHORPY4ISCJN8w+L3M4ykTCkt6CcPli1mcPFFv/r7cO3VfNkf1Cgl+6gXd7LyOTOV0
yFfZ8/8pG0H6QVAe8gIACHEbmN6LsjdqZ+gFBwbZQwENn7FN6EE1LD+huAaefty2U+6F9tjm95Zo
l+Fug7+jNoZGWc3+iJ7hz3SH7biPMRa49n2OlgAacT2FkRX2g82ymTVb1tYuEh23H6LIZTJoOjhg
MG5ajzKfsOkfkHCeD0sI/O8GNA2WwPAdv9jvPabpwSi/erHy/r0YI7hTi40L5+5grazVYAun2oyx
HuN4myUfcwU2btRn5TrM7KeBS5NAdunJE6dLnZclwye7K3KX1neo+vMFFdBKeQ1KMXZ9jsPxeR4n
HxzG+c1UgVMBKsSxZ6RSscTLnCQs54u1yvTtev/sQIMIKWiu6oZZn497lMnsL5rYNfpnrRohLoU1
zUKj2JD38Z7LmSxe8YNk8k4Y6q+u7nRcrPOMsf1N0VNwGvWqcVLi4s1skMCWr8xR7Ckdw8maqBJV
dOGvVz+SOdALkUbMQbRjmkD6l8DnYV+s5cxAtCNQBUp+o5kR6j6DVqPwetj+oOEySH1Xc6b9L6LP
An6uRi0BIrvVcDQeQEIsapSKG53/fQaVPHjC7L5nRlpv0QuabdllFB5V5xzxRMO/E9Lua2C1v3IO
PNg8bIyFCZa7KtemIB+SUZ5b3Wim6biZXMWYX5VAPsXz0M7IDUfam11zG2FpIMzuREYdY5QEmKNS
+pqrxqjE7qHvF+7WisDMYMras3wazTDaJp3RSUYF1PM+ZuY/b+HrMYZwpin2bEEjCLwVt8G5aCv8
YBwXoWQ12dajZvTNBuiuQi4QJwZQNHnLg2ccHzG2yHUGexUM2Yje+DvqRJO+uLOqW1IJH3D/fwWJ
uQjKBBgiICBS0cdeeKsopi2v/G2qCkLuVYoW9DWAK91wsXeD9uPvV/xSNWc7HITfYEZqO6caMC/z
5C3gZG8UYiFiu5dFv9DqxB312dUg+cofzsxiuYDAj/Nh1KiMH+w8oZTqaL5CIpYXMJEa/TIFyFLa
VTOui2fN7hlZZIiy9bE48tO+CpNQcCJwuO50Qk4aOBVJoSQmdQP4NzrGHDp+JEtkhi3SxIdivk/X
hbOOTatCAnxz66hIM0L6m34tpgTYUKNOoYXaAy/jlOTDF2i6DENNqZde/qbvMMe9NbgoIelzCjo/
cqgf8+dxCvZoANBtcP6TQVeXs0TgAF55xgXGpIOId/j0tCJlLwtZTzk7wQhpV+c8MbNifpAwWP3R
w90TNIgx6LLudL7yvAWbSQIknANFQBfX3ZBUZ1qU5VlThH0bsd4fPXanf72xpD5u35nM19R0zPXg
YHmQRHVw4J7k8hUrglO2dF/nBCwfIvBN1iI5GFPwN5/ZCBF/w4SYqyPzdiWWmdF5V4sGj8u/3pR5
odlytwZvXnLosc5BK8T69WC6AXNejSHsy2pVcVujXc7Pmytz7rejAWZbpfWNCj4EpY3ySK1ccncr
8/nTuSnZmvu2RSkPIwYgjYwYZVXTJliSYI7XZj08/xeFda6xJQcehsQTlTuaxG+HaSOPKBMCLs9r
+Wq7Z+YIs0/cgd4S8ajda5xR6gXQLla1BKCC3obnqd190hJEAox3w47Wy+NiWhsRnFk734f52KV+
hIMa87jA5plGT1ddTYLbOzA+gV6EzwLaetoUhY2/+H25PrVgzRuIf8ORYUlhNnI68AjLnu6tejRV
2VoAJyID5gUDHZONVTKiNolZewkcH47eynsBnjs0mLeoNp473FNtGa2VFd5a0533V/R4oBktN8SU
BeTmOaRXE5PZgFCt087TYz4dIJgdsvxnqp7a6udL881k+dXfZGOzMja7hEFiUb91PzDDYoCY8qr3
Pf5SmOPwxIJzU0M3FVS7m4U4oKZ90+wzV6WVEUpK0fzNFatXnJ1FDYzfGnJf2PeCjQRDlksJd5KZ
+6+MhVTzIBzjHFIorXSpiaUBbBOYBp1aFOkCzCGdeeQsLt5Y2bDA8tbbTNA5YmAuH0VGfW+ZFfji
XGj8B5jbXNyQYWLJi6BdLyjJ6B9T3cIQdmV6siJ8GxhWjkzptwAxHoXiKj6e/i7PpQpo2JXUdxqt
Ehft0uj+LCBK6vVda8YNW++nnTXWtaLsgKZjjCRQd03tnzv6OtfrH/RGGMnDDpK/p1nkC3tnKTwE
WTUYKoReVKvUMrYx3ZgN4zhdAR6HZHh3HukOeuPjRfvnwtoZwrxGmV+7ctcP/yyxEVLv91eYoVSp
KKtY8bzx7/xzkEEyGChYWqDWXESy1Pa7iD5F6yHRUggHML3NfJyMVEqCMYlQhMrTSpzsrWuSt9bb
lIJOy+QqStaEFT+FdlML+2LKXzwsbZm5AncSsYsnV4LLnAnAGy086a5Go9DoOZhyGxlcWqzvOknD
IyouQs7/YqRD0A19YCqgRtc72XsN96SwR3JA/kCi7GWDLDNbynny3+XO3iTMxk8vEW7UxJGUMTEU
Mz8T7cPUAaDY9ftk2O9PdSF5qd6NBP6LSo7eSO2Z0J970TNOqLi7eOX1fKHAqoB27Fe+0dDAhjo1
MWqEsZtFgwxmORCy647l9fa3FXws/2l51FV/3mUMT6+D78Ceed202qdkjLv9j11trH4Jn8tiX5uz
/ijTDQdDnagidagBNqjT1OhEaxbKOe5dsBMabSpzO+1bU7cK6rE6ONsZwA04MRe3IIIyAbZmEWim
BYcZ6MWytLos1LjAwtacmFAbg62FmuVNPY4klPV1Ri55bkl/dJCJpzw9c49TQNsbbuFFd89zF89+
cDEftxB2mi42DuEijrpBVEuBcYfSLwuvvUtnHzCDDgtqA4JbhGK+Wy5LxiBHUgKa3GK+AUCFZOVY
PssgJ14oIMHr8HTFtmxjiSCyx4T+4iZZG6bkzyfwQZOAREUi+v/h33PrKJe+civPO9EuFyb29cF+
+wg7+BqJJzAnzcFsoxuXWN8pfZ1gLdtmCROh8Bdpzriid6DJf3T8ApIEOcX2tji1RV96C86Sl1sx
RxsNa3nZhQuxP4zwzE677axxPdnQiMuqQpB2wQUCM90f+A9sHqXYCcq/bwg55WUnnNV6u4xuw8eD
qV5VuaEq8/6GtAfZVDRq5lGKqNSegaMS7bT+mbptC8IWR0T2naqA4Jf5GlymFtTpf6Wgsz5rtKzv
9Yr+9JqGRe6XUpcxf1vlBbOF/4wantAPzLxIgx+aLJO7Ilws9Iye9ZPyAWnHgjVopFxdiubr0snz
ICtftVbZBNlSlXmWq6y6MekcwP1CxZGfnB4J79yMHEswf2WuZtKjAhTI44PFl7RtWAWmWT+XspcD
aH8vMleEpGKffP/CLmg+LsSqTrex5933hF/HrV8G+Mwaiz6aoxCOucRy/Dbzl6EaDiNmtLpaf6gi
SueX34V29JMyCT5AT3fwPNcCV+oLxzciI569kvBM+dMzpfXm6kHEuI2gJIsB3cK8YVbkGDfWOZ5D
UL627YPpULQltqDJ+UPAq8jZk1EXjZTGCe94fdY3kCdgHkYkRkKmW6z3UBVPMsqAxVRRNoo9rv8G
yRPMLbftNHLQBh3CRm3fYVErtL5avq/OknsQMFgxDVl4FoVYc/SdZElgm/T95dbxVIa6npnxRder
u8AQxTIrRCbE6PX/MHEH5TqJbe6BS7ZH/rkD+O7cYMfX4lDArNpjrOfZ9Wc8fG7WSNW0yZpyKvdM
O0rgyxo7W1om1FJAzICRJld+vKp18rJCxjfCGXFLoeIY5Cg4aun6IHYTMYiucfcnjLlsdpnn/GiI
J0iZkKVYRzYmfZYCyM3J4yAAuvl5DloGyTG8cFYDXGD6GFC0NfaT1yNCPAd1ZvPVlxkEQozWIDjE
P/C6HHNkvEW11eMYSaL9x6mNofdkqX9Le+x2DA9Hki4b7drC9mIBkZ00D5NMGLRFY/8J3rGLkiU/
LWWK7abRgSRf8G/X2rlbkXSGp7Kii3PmWnX9AJPnejl2QHJTDsGIMy55IT0UanTZ6eSaZw9XM2Tg
sdjFQN2JjVsM/t5PO9LrLUGY1C6jZT0D9s3684JuIdMK3GJibFYdtoczC7hTCXt63m66vm5OIz/b
soqzcp3maTC+Ux1gA/5gCvIESKBScIauvb+tuadSdr6ux8NiBNBWrnIu3RptH0fMEQzkwm35N7uo
PuoCzxbosZMPOhgJDw2SPFo8f1y7Nx09KBbXcGtJZ7/KpfJiWwGnsHOno3w6ogVTPLEBTCKdORVG
LMOwvc2vM/IuNqjQ1FjvSIO3z0TSyER3JlHhmClzNbPq+HD7rW8csT/9DC3ofFh9Nfvh9s/E6PNG
+maZaHs7NMeI9bwdb9Ew0wSvI33GUH08grJ8nITvqjPNkmL9LgFUmNGK1oRQ0rAutBzs5XRRAdT/
iL/Xc6sdWu70VUkUGAWBPLCLbW+HT9F3lWa0nE9WHUZ4sicMVcD9Uei7lpyJKTeMB2rkqtxvyudI
8zq3aoLPiouuGkjhQZ7BL1lYPjRxGfdwT6Fkm7HjIpeSEWjhWwJ3z0JEo8OdiQvsEsKewGE4s+na
9GKJjot3d/ckf6+0dcFhIvyXHlo6i0Q2mYSLsgDpwOxywRA53po1A7xELyPJMq9qba5bfh3aRzug
6tgm7J1sXjC6zSxbYTk/3u4EYkoqC/eUcAvj/+FulKb0VEBbnYQyu9LZl0UftqMMA++woUt9OqCD
s/P9mmjkqLtRkdzQm4FsFtNR/uorUUtoSTPOMsmir8uXdMknDBONuDUoRJx2QAAUxwvNP40OFX95
WLktqNLxH8llu2hirRqRz9tp/qdqVmEkc96xOD0KL5rvaJFdWOggS6bpzO6D50dAdB/styYMvlvt
YefeaZTzRA2JV2K1I8iNDeB8bqsn4Buv+u1HeDuPtuC4eY9C6vcgLfXN/yWp4XxCPKl0YhHJUFnI
ELTtF0vK2r78hSqlTVHZkcgwyGxkOQ2VsAyxC9SRSZvT93wTWwwsecNnkEoRv7a7exxQ95k8urzt
rasfuoXp6MamSf++XWoJEuEU782ERoNp0MSx4woaLKaE4onRNnKmsRiE0mqyd8OlO09lKr8u5Qli
+wVgzpL6pWLmzESCrFA1QZ8otIypNoixNLlzh3k9u4gZ+mUPEfEqp4BZVAzI6d4vdmBiT2WQ6K21
8UTaB1KzWAHI1ZUZH90CT2m804WuiOCZ2XmJD7oBnBr4CXhoHAaI/8vjT+6p0f3UMLezJCvrTSvf
qjVSwoirKKZcYnkctDIj5RSJIMNOPWruixdBDMvBORNf5MIXcXxFNVS6k//hbfeIJbO1hPNJcfQZ
bDHpznj7w2zEdQ7Nu6pWvBo8zuCXl7IIFUk1nzxcq9k9u0+CTLisEvKNJz6R744z4+ql8CA2qI1r
du9noBe5SQ85yI3Hdvq81OYB7IElPNY2ugiVxzaFqW/OB6fI22NIM0llNyzBrhmChYM76/XMTPlU
i7CCjOwokIPogTE1j0sjzma1lnm7O4aDqCKJHBfVKojRvtNjHsQ6Vn0mGCSEs9eqyToj5jzcRHYF
Tu/fhzNbvamhJ+A+hrsF/3NttApJGzQzkbWoK6Fn7xNBdMbpXobAZCbG4I3AuwnKAsbpe6l3+cSp
wU/Ygb/cW6pxadDsuLLVe4ywiW1uusF/Wf7g/58FJrZwnJjyGB/S84ClAgtm1Mhf0ItqREtzFGqq
4fN9I5+GUxWb+rhitOlQ2pFpTyuD87T+GU4u+04h6YHVKQlHt7p/dVWDrPOIXXPH1gTy30D/Ysp4
q0drgwHTB7oCk0jSYZ6s7XUuFqeYTV9T7SPR99/vJMS2rSQcEiXwmlATWy0fexu8rv7Yeq9jbEHm
IQEWOrxG+mEyED/hvEgoQc9+6ERIYwx15a265r4j9atlDi2YjxvU8oG4Szi5tq2ZE63K2YrbfRLX
tY/reNdFplkMRGILcAg6eycRhJa5S2tYAqZ02mpVZe6frpbs02lvX2A/nv+c1huEbPhwKcjRe+E3
1fJfoz2wHif/8V7bBrhdl7T1FVxzJcLZ+XqJfKmkWrOTM4edDzfkNBIqMzszfzbMGg5H9lLWw54E
NxkTBjEDvkOgrqNEIlbcmZMEN2vjboSz9GmLLgjPGI1ACFw9yz0QlhQMxFw8HCS8pPlp/XWUrEAN
STinRiikbJwYyIYPl6IUPKCEnYUxKPHI4C0yTF4Xd06qFVmMJ3/pUlmyQtSphoOnXpSD36aAYkmj
sQDERSmuhrkk3UQ1vTSWAQqWDurI63kd2upx99QKSR42UI+qzsMdOKfGu/XQ+qW/np2tEmfyDL0M
moVdbhGXMSUs5w/piAnd9Hux5r0FX8GYPn1KObHYs8yMy+pLfp6Hvtp6QLs/rmCQikYp3u/JCdkd
SigDhNcEfDrPY5PUow6YhvaJd8mxxZpRb9dvyKBoHVbcagVaHiVXCtKqZmW1iMw9vY4O8fYH0Lt3
NzOa1sUxo1uiaF1rg8B3CKHQS6Uf3xgO7FTewL1Zf8sCWbWYHqYz2Y7Nl8XKItRnKpTNynI5+dRS
zalixC4+sRjF+Dsb/EJMlulPtKOmPN6ObtpyAHMQx3nORtIGYnfWdCUm90P8xDNXFWgSTDW/V5/t
mNV0+wP/PG4dTeywMKJAhS9JdLl2pZu4JdxYF+T836AVMhGMN1g6uvaz8MkbgSKj7CU/oaHsXxvw
Kak0Gn/YHbMzKbppgM8c9WPJYCV2yYtxH+g4S2iJS8s7y/Kc3mVmHk0Kmgz6cd4B7sXpwtaScsi7
E3iH9MXt7KGVvFQVDKTny7XvERuo0MquGQ3XNwTBZlSgFTjsk6q9eg/B3XPa3t8FhVM9kALguZtE
mCdP6WzL6bpEEWbWyuE+hf4AgfxtqAJjNnEeW9fLtjdRolUIIcTImS9S2r8YZr05+ElDAjbQb93/
Usy6fUP2omXR4q3QHkjI9Ew1Jdtg4gj3C+V/MRU8vBuI0JL01KOYgwixw++3q/5KjNEWHl78kXsX
7XXHF/PrUkbFGlZmL08xtOBwzwSg1RHTZEipOLmr1aKj6TUBkz9dU4tAMc86t33h3jMm938T4hHW
a/q/7FpopuBnrxoP008GogtK4Etq09n7IeyauyE3WkSeqLukkfnPfUt18JbFcIxnVnTG4vGYXjUO
cFDSYesp4Gjdp9hN8g/AUSQMQqlAy2vEijDckwspbSMTnar+QK1UrrF7uuPznjzAG5pzoeyD1hh6
gmilYPSKrk5Xt+q2PDT6kl4H+uV7zkgIQ7Yg+j/bI+ZYCwWR3FSZQLbpEgfVApMXP4WC0eaMsMoI
wZdsbgjnMZsKMd2jcP7AEv1XSMi+IehkxjzQ1XaC+EBel/Gb+Do9Hh5K+a2oo/sjIwcXZXT7P6nz
Gc+bQeVe0DviXy1WVv4uzdmh+dGVboIUXBv4HXQpaZD2sJQ39JPSH6xJxYqCUKw4kZ1xug7uwLsx
RSlNTgsU5aZi3Ie6+46QM4IE6pnH9p6pow5/YLIwZNlXZAMMZEBYy5u0H2ICUjzKXO37ohsLRYc1
H/J0pUT8JeiYuTLuAFotdzxEqUIyyCYH/UC3+eaEzkWtXD70huAuq6Ae3yEvDhz6nN9ZVLXo9Bqw
IG8d9D84iqAq7tGY/r6ExuP1qA71KLIeXFtJSZNt7kKo8Sb3zbbGWhGAlFTLNPVbDrUXg1h4UiCp
l+BzgXKD+mqsGFO/b1uOO2C3H9MPVcx1E3g5bNm03XaeOeY0Z/uWGP/XpEbVV36uIFNSHRwfE3bN
eEV8WUc7yImP+Fn4J+OzTiN7u9BrfZvr5ndKRnJqFQ+oycRw4QhcBNNaaw1eRKOmnKSpE1BHBrJY
ItNnVtA8oWA+jvpRsBTDEenD/8j0xX8E8sVGnQB8yWz+pfVBH3VL69xWE+9YKo0zv2MdxaWIvOBA
HZoKPYx/8tfybdMku/UeXRuE13fMUYIo+wD2r0zqLDfmB4Y7+Eb2mySmVjZorsRsMFTFjSsYCql7
xvTgCVZwTyp3xP26X3TsYomyX1R4ouR31MdYTungqXCciO/w5rOfpoyIU40T40Wg7ffOO5HqR+7R
oVpRaWIzDQjjv8rcp98u2q0R487NcKHEl08QSlmf3YsXhWeZnX3tO+FxKilbcwBSiYF0MnxUH648
iYjlFbkGtm1//Z0w0aMP/gDtNt/O5g47ZztS1jr0OucELuB5mui/nBRoa7FdPpmLgJUDX5aIRtPe
dYVOL9VTXTLjus43E/X+iMCoMfrUID+WrRkH4A10oSByuzhvUXQXCWO45peyMtHvu96qEOsAAVoi
+W1KgSLGiVnbLkEP8zEBPGf2H+f7mhcZDLgCrKASxgrtZ+tcK76Z82rterQT3XPKstftwziPWu6T
ayX1hPOeSS/+XSIY25OYfz6URCeMLn6i4B/HV/q8W/F2pfPIKU9XmkVqF809182AfJIoVP8oV/jj
RPE3ckHuLTcOahGv4gh/j6NiLsFBqcR/gQ3MnS8NnX/U6AZn8ggNO6sFKU2FiCik2E3m7ZFxUeI5
M3wX8Y1dMZkHFQ5E/keVNERMYsKKgB3cxqfJmB/ownZR3nYB0ATeVt7U7kV7Q208JHqxNTY/0nbg
S4QBg5IOesxaKLmkubTsvjU4qLzQkHVDY0WVqaT+LuEuNU7CCeLr5z9ay0fbuBMvzeypQ7x9c8FF
1FG32ASv3+EfKWJZxSNpUAMxozLfZ5fiHgB8y8qT7HctXFm5hH4PeXwF/z9bbK73DRqvstrH9lZm
VqlgIqg5lkeTqc5KN4SMU928Pe/ASdVROfxU0EtLNOT3MI9+eTH7FTUExEMlfMycyKdhjgqCAiT+
5dpoAHe8e2UcFGnbypzi0lqefY9UNIeG7FGzk7xmz+jhcRKuiWJt09gzOXwirs0o7eV+c8kZb81N
QMzzbVRlonR0n/ihSrjZc1/ZqK68BPlr7To5ljElvBb71SEITGPXtO2WAsF/qI0if5NVPJ6sTD5M
NlX3Mf9MS3PAeV5D50M7DHMM5rQB+oYLPF61WPPKw1znriI6AMGCEEceLw4ENTsDArW13l8HogCX
B+HqLlMTLTy6qO9ibZs5AdvICgN9l1Avyew9xRGPIytge9jxZ6MzD6ehFXZeuXdVUnJaO4RmP93p
B3xY4z249/kxWrfJE5Ablrn0i8WUj9kHqY833hbpFKFWUmt36aOy9MtlvqRkTXmBYXRke9wC6h77
MH3z1h7qDWDaGhLJ/R1xDV4gKt4bobu77E9rkQ2fCQJ9ri8KSXjuStdwfxdUAB2/QanipSJlMyQw
gIAuRTiyXXxxutxPhgfn2dnbyaWz8fKdNFqsabg/zY48BQUgOrWaotanC6FlpHl9sd8o2TZxEQSo
EZkCmywZrVAhUWU1S9rpWDtbooDrGcVn+lAvjSRaCvazJQRvHvpjUnj25d7sUTvxAR7ukf50JQJ5
xCebzz7E1pvNensuakTicQcFOasZehfMgHQpAf4HV/5CyZXTnzWp0wfuFNhaJ1oH1ZPJMWxAWQY3
Z9YRORa7fWuv8da+aNY1cwLyxjGSQ5zlqtmSw/zf9vU4CaZFWBV9Xu1R8mhMH6GO9BBEu+NnxGek
SBZnA6gtbE9wqGjBdYOtz6gMu/DDURJmSig4fSREWA8p3ZzQFBkjXeKsXdI9+s9x/OsRR2BjQnQk
+g4nAKh8L9RTCpb9srqIZ/CerHIM0K/YrII/uLuLAVIBUBIJ+cMeqE2dkwwtTNm39g9ZX1TuYC9w
S24b5/3Brm7DT4+SnWU60ERi5oea93UoOAp2bX1qxFwwdspQ/wtjPrWftoag3PR62jX6Oy0L7xSF
uekR8CRgqhpvUgyhvMtZLT/t9VwVf4iVjESJg4JXvo5LR22V9S86HwaqdtDVVKhlzDCpMSaSCWGw
762s8cU44vRE6c+rh4UmGdrCsX++jimOgYSz4DqOAcMqAfe86cGIUKgag/eWgYPqqoqzpMPzYShB
sm/SO8d1cSBKHfqUjN5zzmm3ozsKolzlEw7juD+m2S10oebUVQ6wEjM5hQGIYwYBWoeNRRu0sHHC
onp+3o/kGtrLTfe3h5YjvuQ0kcp2TR8KCAz39BSN1Zlu4YhLl0Pq2dH091FDhU8n3IZ2PgRbS8bQ
wcpIMYIk66ac6SPcUZN/u5JMZYIp4GpMS0WKXb6Z0IdPeonbibQJDjqSnZYR/FSIHw1A5DrjU5ek
DWiJvY0kj7B2gK4PY7L7MRUWs+wotCtnM5EMttFeYJE65aW+n9NHsWTGc85pQYc/bGD0akG0lV+j
IStUj6dvzKg69Vg8dsX4LFuohnkjblaf4eZbvA2OVwxrxrSo9VdhTXgkJKnzQ9g67lUUIcL9cQFw
GV5ZOCo4BuvZkL1lMfhjxEahROfI7KzFAAL9+O6s+m+571WP8zz60RD687b1KpF1dANCj45CMrkd
u0VMzpAnrN6PE/P0jj/LaQAcMddVJlwzN7HfjAg18NkWt5MqeIR/PJxwDIyBsICw92MBfyh0SldW
aknO+UWycZ1BMGd8nP1pOS2JMUg8jGoY+OF2u7fRa5Naf7w3KT8vhtgnkmZAeRofp+GmndH4VHtx
PG64m8CsnHEVUU3SDKFI78yNHKiDGuscjHazQ06uOVi5CDItNoOvHEJOZWydJlDdu/LIAkd05LXN
/ENAnYx1Gl2BSzM1+zN1g22u/Iq8Qyr6KrDyFVPxzEs0np8NFX44ATtI6r5k/8mfLcbLrhdOxEiQ
jDX6LamZECKa7V3rSIxJKykRhKzj8Ix/dkJRWM9Wxwkjlb3fECblEdwotgv4pCdSu7g01CSrN5tK
QD2P2ZCH9ilAVvxI0oNYEJ1ouNviwraBuRWdY1JPL/zvjb/m1YfvgcavBgorpLF5aNrQbEtBpO17
KkXVxqPfwuYXdSsZzolupKqig8CUQ+e9/B0OUk53foo461HalQV+FFCIuxmSfyWNnvsay+LvdyTj
iykIo951ihiP2Kq6X8M+JvBWt2JTQCYv6EcKi8MPgqURXZ24FRCN8hJple0RiHNeIO7NbtxuznF8
Bkrw5278GnjR0RrIy78iLa0ZPxlLmitK3rk41LY7Rma58wKNvKWs3T1pWqHz4pBpq46KBUxiWtnn
bLpQDLPBNFGzXHF7Jp2K9LlZgEoPMjBpSi2SV7Go27XqinN85U1eJlJeUjEL1K+yzUQqfx2k68k+
8d86VyyWslYytX1Z3GQLMRySW1hkVzh4ZLHXt+DA394mECQ/veK0nzo6Y7/NDXYA0uTgBROxfwIn
RqGz4filGrTmFuf6lQP0mtFTgnpz19Yd3aFBfn9EpcuSixdci73foqNKBBAAUJtLiz5348FRo87j
sSzVzeIl3RFePn7C4LJYjv4YaAd3I/5ublNHUOySu7a3JOCCqgmtsY4U2W7U0awWc22TDA7SkT7R
5NdSRpWZF2E5LQR5SBO1H3AvXjX04qrRsJt4MJ3yu0xO/ZMJCTiekPoChkJIIKmUIamC1wG0d2tg
rVrb1UdyZfjFaPdLrI8tVMj6xx5z7X2ktOeYl8zyE1pAXj5sCTNC7S4nqItq6D6YpwiJqVhnYDYT
EXMkGJeiQrkRP2jKW/fRM5zCgOt3tVhYpViEK1ckZc1eoqNedW7Gf5dkk2aI+YCxd769fV5sCyZN
t8AE6w/pUWPbzF6WrJhQMc9+8gITGCHfdMu4VZuXKBr1ijqgVvsjFthl+9YkGoRYvABiucQquUW1
rth0392DndIG2AhPb7cmxOgfrSksf1YSsfH6G8bfz33+IlIY4WM9eGNjnO36nE0u9UF/xFJT6/j9
Toj4XIUdvR01MoP3nsymcEIYP53rwcIQ2lr3HOfq8eDgYZnqmcHBggdY0cpFVkSJqsIkk0bP/0EB
IE/uaKLBxe+OD+k4a5oLKL848+rmQaJBtjvQ9AfacAy1AtZDlD18pZ6Xsw6aYTREPqGI2Da9kTwV
s7nzijjSW5JImvNkt2ugQIFBLCtEb2cWG+MHrJGB13xJzqiyq+PgHSQnvm4lJrfOFnr0HBwGXFvk
1HpbEqd9G3sR46Erupp43GFI1AB5++SLPKfNVKvXwMk4w/hBI1KnU0gFDhqKpPee4r/DOuDNaCBP
fV4zw2tg8BQ+HzM0m4hlGuwcFMqWg36H5YFrJL0INoSu7wns9dCe9T1tOAUczBRrPhrQ8rL7Siu5
d70yZFxWpoidBfD/t7I6BkviBYXuISz3cJDONsGd9/vjfypw6EeTE89JCIX2m/rh/6ur2vXdVW49
GZ8fFO+K0TXdNgkoaGZWvUczguMnyMPCZNbsHkcflcbwsUQCZ5wQIxaU+9SrruD2ssCpgDwGIQlZ
iSDMNbNTYG+8YbVSlvbfeXbQzlAY1oRe4q+P+3vHoF8Ks4vokCawT/FkQXKPtJHl4IPKEyr+lOiI
ZCC2J36xa0oQg9AnNoJGGl5T2RmFhAWWUhChZ8/+WLNEwChq7C1qyWElroq4GZqOKmjPuGtQu3j2
bIT8zjs0cKR5tTPh+/fEbfrj0H4BaNaSa78DeH1nGs09T1teTul/Vcvj3Pcvb3K/N+OUrwiuj/hH
pg00TsW81sl/qiXC8F2DE3bkXqflKR7vNfBIF4HJmXlP4YUVhClThGOR039S4iKMIJ0nRoT7E3HL
fzjAIKoL/JLxU4FXjtGt6rtxjR2WYXqWZ+SBW0DFHKD4RlYcU/SE45QHTF282YctmvlmVRSLlcbp
cqGzLkrfBYofXzlPMdRY8N2GoxNPuSClNdYi+4n7t1DNtZLh8IS8nB0BmepyAQYwfkZWDx+VpHOi
xKHRTMmZ05RwUw254vgtRid58SSiiza+jClX3NtD6v4qrS1Sf7L+rJS6/nTDn995bPU5xr6UuulS
CMFTASiOFRQbe6dBcZ2ceiJ3UQtvpAs9QlJCwSTb3Lm5ePkZn5W8SWWCfPTrBywAagkULI8psZtF
olD02aWPU37ZAHISuAARSY1AynUP96oqWye61YQXTfFwIEjn3tWbLluESH0jG59bZqfgfNawJaU4
fTrdLVzrGkGHmfYvJBB2jl++EvejP1Hd76lwybVBU6QM4zxtkEgoEMyuV+ITTxx45cds47A+1jCE
FrjOwhZj2L9aCqzRihUYQRcrGA/gO+KNGgmZOPaZkyexEgZnnY8PSGxcnP1/UBZSQ2EsoWS+uwEM
w9gm4BCdL7jJ4BZHvxnRRQQhei1PZJCxlJD2yIMhnmQkYpVQROHbjtXL3wgufM3OTPT3xBVYRbs1
xaIAlKnTpg0e7/5C28VcXRQWzSWOBMy4hH3Wxuk3PgXWbWV/3wpn0jlM0E/PU19DRnZHvsWPJneL
zwnY2kSltM5uvIZQpVvLqqC4I7amL6+Wfr0oblNH98eBYvjve563iUnih3RT3RwuuBeIo2zw+l34
NeXM5lSGHLnva7/t3p1tn23r5+jjHQwb5HJBUri7eQJPWLB5vFt7mJJKcTGjj5uZOS1PJOV75ZgN
ebsoMi/2/jWCAWRbJrMHAiL/H3O/MR7D7gsPowa2wXxi18LTNhfuFJefsDMiSgp1GmpdAkiC73WP
YXrDyN0Uonl6c+/BC4+q0YMpZqVT9dBsFh/e54jxBtb8xIQnJNskWtmASmHCgyGK2FDJadTWDUpW
m4pS5or1M+iL6RhNtNlAru8EzkIZ66DrsKjOLumn8Pw/GV8cjrxfmifPOCPcEVleQEX/Pnt3c1Sf
R8dMGyK3UdRGxeEBc33d2yD/2bLeTz56p+30ryeUHo3BMuCSTCkFLnhhtJbf4NKNARTodLdo06L5
qXmMzpfwGhCt4EacnNB+2WixoLi7gGejl+qM/bYOzNloL6qpju/pWxaxQo/7NWa2u6/GhlE2wBI8
N1BJZcVjhmqGJ/3pG26fQ1z6FcqCH+ICGG4Y/tavZ5eWOgtZUVNJpJzqhZnlSREAOJxfFV86uy26
DLNGIg0VFgZqv41HIDfHTGiHvSFLcX/BAa2mvLLOKaYNV+Db07rb0TbW4KsqrJ7Nry7+SwfcPUey
NLawhfx105bsNExSjVA4oEpq7muXbZRAOO4ib/P6tclygEL1l9OMbEREeqC2gXotuwk1OrxWioYv
lpMg2M+BKSb75VslsgSYSvp+1Bgqd2l3P6F34QukDOaipSQpbAPqnKx0poYu6pU9NZTCmpYdZRDu
ZCqbqw84Zx/eoeXYU4rbLd80/uyyaH7QFj8pOK0uKnXwsFohoJvrbQLD4VBzCnQhWa3CAf71AzTH
dXWCiL8tUe0mBJmWrhdFS3cBG25/fbjloDurRe0CEe8NGpUOutPH7+v2ayR0DPLNykkZnRINGHpT
1ZYmJQg2nXkILg1JuaA0WaTGCUKFFpWTINVu9yt7dLT3WiYYAy6gJndpsUCe/WozyitKBLp0iaiA
ByfNtv8JSIhI2m/xqG6PQUQnZhC4dJYCHcj0drRlZ8IjQCqXbgay84tsqif3aAUc12NFcgQmsnO8
mcIUW4IIwkVFkDHOBYzNU9qQXY1o2XgaOjaCyO372hZaLR1Qf5PFxkFeSi6UNt8rVyMbquXW5QA3
//0+t0eBSxx0XEC4FmnD0LQkiNLhcUFzYMAMJw9aEqm0V8huI6AAt1J1/i0BNw6XZDlgRdCMew48
Z79B9U2k/cQYF7tISx4X2rNoIVXsH+TuJ2hb5MYcshhRqkmDnGoJ+pQdRUzebK2gfoeNUtjE+QJb
5yfFx9Lm2efabjVcZHCAhJObYoOnupoW8gHSKedEdT6pa5qbr+2BfZVAaV6MwvTHEM2t+ycuHjKt
I/1792X6v7BY+n803tpJYxjAwT0lLcTolqhafddLkx2Dennrpcuix0hiUej23Nx8bKpQiu1gBDEZ
mp7vLd5eU06nXyV8RSsEtMjR1CNY9WadrGbv6/BCIDlAq7j34eiM0PsCO3wRiOsSHjOmn9sQTg0p
CpVBrAkzgvrXxwbUbwyKnZKB0bVU/6kREh+fxxl5c4E2dLGkPz3Ks4HQVJeeqJeXOOpCUpDUXHny
XLw4bHo8XBL1xQ7YgyKXr9aKSkGRjr0WHgkD9lMPC9AvjrDx3nlw94fKYYZcFVao/FwngYrAH1Rb
kcz8v1kANd1h/JUOlG0sRIlyahEYLV94C91XcU5UcDSmlewkkEJI+K1VQpdWWIFPAepZI8Z6h7Cc
EQSXe4SibU4yL0afgR8zwXjMXlpUJk1JlMP2KThD1zpvTLR8OjuNjsfPsnsC0ykEDGyKv7mvIFy0
+Eb6xANeAgtNrqT4vDakUjqOAqZn/2LhN4tevbigkLGagrhCJCRCUSotQB2J5m/6poHZXLfHUQih
eDTUgDADT/EoDkFti9ZV0lIxhCCoZes6nCiQtSQj/4QhOsPe+1011yD/c04J7fvO+jS6+9mklR+2
u1unsg0J5xS7qwB8LVj4M3RBeP4clMYZxNXha/vFy7oF3aJXvUM7UQ9OwnC3c4XUt8KU8bTD7FQs
Uq71GrQcV3aJxQQqQ2HY7WqvRbqLJ2c1z0Km2BJBqrJg85T7DsTIibYFw5nZoH+P1vvxa27J0StO
9FRzyZv8lG0oY/OP4xUTQHn28vl3OMWcywoVTAUiii7ZFoxdCt8qYaBSmkh8ZDWx/aLo9bt1dHGy
je/AKRAnlpdiyhQz7st8kJxhrq6ibruSXIgn4S0eR14tH92ACLC7OChiyl85AcAZttMICiztyrzJ
CkdShuYdjkKAjpJC6WOCa0rCxknBZodbcUESyh6PiDfVaU9NfDoTo0b1z3Y7qCI44Rjy0ggsvBhT
5iuqPBvpnY8zYVW81ubEHHPuXqr18aoVaTrU9aQ/7dqDTGxwwT1SfOuxpwLx2uzuVbRvNIsAmTbh
oO2gGdorXIXyCOSTl12GWJLsKdGpT0Ht0DK+rsO1UUT+LnqpeZgOC/2xSBaAzXppk1HMCdQLFsFY
A4NMvS9vgpmobd34PBip7A0i1S+A805TkQd7vQQrST0T9or9TRp7q254tw24eYAqO255f63/MW2E
VxV1OGQl237Ee46TeHgIT7sAZdO1EoECGI9exeA+JU6Rd4ZiGKaP/MAQbpNZ3JFq1Z8UhmfdPGZH
B7BqLyeBAFXVcYz9x1GsQHJzB/pNjv+wwGcwirUewHDrEW7F0YviWvwbWDIDtplDREdvW0UsOCEr
/O1ILF3c7Aas5Qt4+7LXUgp9oXjyMQv179Ky6BaiH1S/fA4PXCh5U2/u0QSkESBNJy8FuBUoKJvB
orUId6LntwyUpw/MkoREtDhRRcisSqOOYN8RJia9LA/IW/xs+NP9rMgpY3zvblAq6tD2VWP+MZjh
ImXJ0qjfShHWFQpUN8ojuLbWTdjJF9km8N3pOupWJqNVFqZ/IW02d6OAOC06uep04qM/fnBpTgwM
S7E7lSiaTf4hScdN8rmx/CkQ10c4nHG3QeBTn6IdY2esagPnDC4uHnRmg8LDoZWgtOZ+h+UtF1Yl
jXCXJ4nLmNvUU3SWhMuLsHJhN4GoTEbOTGTbZTHjGHzoEHeKfbsrBUB9NCqmf/TG/GQgnA0dirYT
ouKPab8CXr3ot75ke6dMNLv35sAKPcLBlWVovE3die0KQ++zgpNaDsWy/6N7c2afNz9e2GplE3hw
gQ8egHiSVvo9/fPTqquoZuaPt9BEzkNdaaGwtKb2g44LRtIM3oltlN7itBSf+5/+LuuqGbxB+kjL
OeSoYJGhqezOTUrqFeqfNjH6mXXlH8/9L2mS5evf0SbbAaTQt1y5JKm/6nNUGddPf9Y48VvhmP76
XxjskqO10GOhRjEgntxR5vEGEyjrgpsJ5CRhqMMR2wMn9ogZevZwXFrEr1OT32Ve0oLLbMfMvuIp
2aoltN+FaxupzSEQu8p8BswfKzGWruBJpUzwMVh2yGDzO/pyrkK+eu4vN/Btvjx139hj00mDgeQ3
MqkMAUD1z0gyFAu8BnYVrQQtnMOnfTDFarXYvI7E4T7XaU+qyA+fM1gOyaLwNgHeH/cglFN2fM68
TSkkAI9zxv/5k/TX8h0saZd+BMfJpxNCNVfhquNz0ZS7OlRRUrmJ6bX/wdJ1EJCjUyCYKQchblAe
McM8PusoC7In9NigcpTPaJlp3uHm1fDsxEy9hfJnOxqPP5G1bn0cfrikoFeDS5emLiUlYS20NH84
owJECkR+paoPbLujvZjDGIs3uxyUf1GWedp59Ekx4K0mKLI5lSKPxdzsn4d4otwx1DqO8wSEw3ip
bUW9JQyMStCy8FhOKWEJXIj6o8eZWyjne1nWHZ5pswMXn3/El0HMxlXBNi1sfkVLoxdpZAuDLs7d
xevbXxXsPlw4eTvFZFcG4UguTrVnNGeInS9caN5Sutc+LrVJadH1ODyFtCSplPV4bZMukZ/o4Lic
w8C+ux/D+cmQtFzngTGcn+eMUGDOObzH6PfHnoPHNfTza77SWm/9kmbGHElKAO5slSMrH9uRY9xK
nM8XXqumydQ7O1D6fYgQI1WOqenfukkv2h9dcHTdPAfBVsDkaNP/eOINCI13T+4P/pzgeSTaampO
tG9cU+Rht5+35wyG8bUu4uO3kK7XBoSN9+uwUhNiSXBqrHX8pT5VRfXRj7LiF1NdClfZxqo4HjRb
4G9NSmCQ1/frmTQ+CeJ0vREzqpOp8BcC0KDSNIDfFwN0v0FN6qBdLlv6ZeCx9zQnYqeLdnX0tD7H
mtz2C4bJ3mqxZA4oPajffVso6KtJTcn5yKvg64uR0sPQsjbrDneMjmvyBtGzJAFaWmR/28esGk9P
zO95Sv/41yeZObsiYfMscfbiSmrxSJ8UxzBFbSJe/j8e20kKhxHNpUj2yvji98ZFszDVEYIfPJn2
QBl3CC8r8mFd9azRkEgAjxnWS6aN1DnC6Fgdao02ffAqaE7tBpd/rFUysFB27+NUFiYjkRvlG9fU
6VHzgnY9y7qLH3Do1RvGnJYj3ZShjsShqgAyKizlL7OrDBvfCdfCaX5rUqE1FFIdWD5usDX7ma3h
3D1RDbsdFPD8b8iVnFGfF81Kh/AtAX3XzJfYkRoMj2TCDRpt/frV/DIYrev/ODG5N5LRuOI5lYFO
4buZPUecg1L3mZTWN7qyA6+/HAgxCYrmmM4cLQIipOMTZtSU1+ojP0WaK5OaXPPq7/m15HIqvbOz
QJ7J87taD+E6KlX2f4kJLTQyvBQg5WmDmE5xc0vCtCWSlqYwDJsjIsgZ6v0dwaQ2alVYKZsW3a7V
VylkAWg+z2BRwOdPEG4vqkh1FCn6WPZNtz7WpyJljEphUXsnynLQG+C3h1ut6bMovt54DxDBnogY
NIgz+8qRxsdVu9qP9LNIak22kneJDBCAbAbOJO9C2Fdx1Pw3OgmY46hNj5X940pUizi3ite1Vpmk
bDEMXfy9SjN5Md8/oMqoNpMUgDDm6TTPtpWkHFvUOoBa3Cm8D8yELwqL33LhNSwU1EHuaZlhib1j
oFFEAmopm+j52GjPPGgyj8HOVKK2W3PfXk223Awn9+r5EYuyzz2idi+Y48vouWCzrl0Qz28xiLkI
hrW0fG3530fV1Yg7wvJGUzFMcVIMWsnaWrL+1I4LZP2mP87D8JVrRdrF7H3icRVvvKwEP+rgEqIk
Wm6uHpakHIOSPgcVFQNTr2YKVT4A+nbtXDLXy6XLu0fDHCd8Y6OauyeAsqzpRspIfyLcaVHE1pj6
hTpj9+X/5qN1EmJj1sau/sw+a+uMR5yrJ+DKIc5YtK3g7G8xtvBowwWPJrkumTiBwu6LBi3HTbta
OyM/fqxPrpBDRTof610ftmlxfj+s2PWkNSs9z1+dPPqXsaXzvZvN3Nx9GiUO3AcCMvwEhgH4Y+el
Mxt6hdTPzWSZAEABCxB6Z9QjQRHkoWXtJX7jVdFRD1GIBOW3ctPCzEcSHqSgyH6J8Y7+a5/YnPgq
aMxkCWirTYyNGoZPDMsJu2WVGjYoRuzw4GocnrCEvBbuDSWGWqry1+OJZCQo/+R8x8UufaZm8OH9
9HvNKawlZTduLOszxIlzhB2hBzyzW4R2e6FCLAgg6P+2uoOo8GcjKzPr5A7qdGuNt0dVwKsP4xeu
OIxJm3Y2RUqGm19QAg6PruOfz/aVilElZliV6X7DYy+SC+qJUIpmjPJ4IC2fx7Arq+B5hcPYrtih
mEZKO0ENXCNV0ytSk6XAgQEdzsWqVH2cG4czuvlIKyM4JMuHJ5Tyez8RdbOpn2E66dHxB9x8QLsi
nSjw0HPVrjpyKCwA/O7aeIa5ATckie7R9QfhAWkN+cP8LqUQPmBU/AqUBuIYzeU9IfykdGOAZmU9
Wd/HpAw5cjjpeDcoG0jlnVqnMQhQF9y6uq4HiGP+s+aVeP2p0qqf1PkImXWI+AcxgDu4V8OYO5yj
3Ti7YOKwJxfvrwtkIL3ffsEjNs3t67dqbFQVCM3AgR4wffBgN39hKDNc8LCW6AKUtIn+DF6n7oFR
hk6HDOnnJSQqWD1qWoB4oNz3hcYR/o9u8XH9Hc1YxQ9Tb+qOHQ1jRBzlthhbtB92HdyUijfD6h5m
7B0Zzjzy5lKzoLBl/RRgIuXaxExbFe9/Nk45wEsBG0wtD2eR1o8ytIw5SW5pwcb8mUd4Lv6egt94
c4fWOZ5i2R4cbvja7pnFaCOhJz7iUJdnUa8dnIpR5H/2r/iEbLC2GI8Oeg5SSMBz5V3QGqtEA5Qi
srk52L+JOGQfpGxFnmiEohhTVpaFaYXlBejyvU4VnuOpNDWFNnrc1umFv1ccRoSDtgRKjEdbRzY8
wyuwdq2AyuGkx73BAOBv7IOhhDFm0KqYk81LjFC3a30hS+MrQvPua7n8Wy42XR0PSPJ4Dy8FPXuo
yW4Mw65QTyIUv2NdnkLbHZoCDBa6I2ZjF+AnQKIqH8qSo34S9SBR3iJvfxIcogLCj9TYTWFi8t54
Lsy9XnMfLLrtM0CbW4C47JaZ9DUHwOgM5rBP4zLkR/CGc6d/ZO69vcAeaelsPn0BlYt/JMnyHhx4
3P25UU2iTz7oeW1SibhR2SxiVLoRjrZ8ytQhUGQ/7z367H5ATjyHuF+YG9n+bM8KAPvlynEyR8Zn
a+Ack9Fdywa3g7Ee6WWQL9HiAFI9ewRK5edhdj4H0QkRsU5BNXZhP6GI3Q4CtJPtC6pklDlPfiy8
A9vJ/m7wQ8WAckuaTwDlLSUjsQn6ZjdrL7vSxpfW2E+P3Hi+0ZHawFyu4Rjn9WBgXRemPGfIaj2x
Iw9zyXegj6r+ufKpt2x4GJk2o3hnbCshJqzEdok7Pj4wh2CPgDO2JUzXtRzxbym5slKcCthotF7S
ZfqhhMYAwD3JGkPhXOrysG6/tKxe4erVF43NB+dZ+GILuREwpHnh12P6SC11q3Qgbo0QEibEtMwR
6thsEUUn36MKazqiShalFVMlcc0TnssKjSfA5+JpiDEHpCdYPbn0ZxyyZvxbFBgDr2jzes8Ty9Nw
viiSM+qy2PSXNPU3v5zC+5sc6ab4Da/nkOnZCkRAoBK8CX+bHi7DiON4igql+Oy1wbcDH4/lDoff
/CB0x6+Ih/M8G4hmvXoiUcLDh2Ytu2fVPE8Kf7P7Th/TyW2vUgKwvRKoxY0doUFQ2226JbJRFMqL
1Vvj4Fg+D/k4GRCilhaiYdy1XNtj3dBN+kSF2ymGxXg7IMctkQqbDY+86rFPJWCsXK9/IZ9pEtfe
1MGmUcMt2hU2yZcvA7YKTNkl55RmnFbWigJWmqk1EUkrTTyUYBKI4WHCWtyJ+eSu1m6XrXckDzYF
BkKy2ujb+TSyDNk+9NfedBFBalQilJQu8v9rqiRH0a5R1LgqfHmGYAfqzErnRaz+zPf0Taoup3Ds
jEbFmopUu4BSbW+pfkBrnxP8Ox4JcSNyZFnxQzyJkMIjcz0a82S+Ftbm0VYZ3G2e/+9fNbBUcD8i
7qs2wxgRDUllI6XTpoFw2XXWk3lyisTHEeTcZlSdwJq/lRn5gKAZzQn/wtVYCcLS/vNsRJO8tpW9
qAXWeS3u9jdJdH38GYwD05tf/MRtR+8Q2cgB2XV3bUl/Ji7g6Iidhp7Ewki5c2VqIrCWVe8se0MJ
lcMFNwDRlssnn08QntAP4FJVzI6SOj51JR79kcLXCqjQUkCGlB9ZlOdBcHuyvwFKUETEtVQeGzzQ
m77EymVwYKFvOiuhtnlvgpngs9fnY6zPdiA4q+S+smNvimONZBLAZF29PaXPK5Ehbrp1fpJ+Elzz
d7/UxBmPTTgQafEWpqOvPR676UPCvlmzvu0xiKyHfUI4o9R0xie9CGYBdLpMWpm7MPrwOBdjPMxB
YpDXqjhtSc1G0p0taj6kmZKV9KcTdRZmJ+MunvvpAd5NSHM2eAmgH/Fc2vQBkdu6fH+r753H7mMl
WCqN9wTKGNzpX2EABLBDShk78X0/zi+1Gf4PIpPhv6hMp+C3996fnbXYtOO9yRQEieXVAi6hHsLh
CMXHde91XXJ5TTX5DyjUHSApJGWosXs7fg4h9YFfxWt/+CWOlp2ipg9yLIv9cC3y9TouKkDHIBOQ
xqP8iwoaCJuosBtjcZBRZRUgJtaOYFyIgdPofO0/EQXXzpDs4rml4blR9INhMVjIc1LIhDat75S/
yrTtf95VX1J+NHeYlWB7BNC61KXbGVY7yTiOTZqxdaPv7osRwhWySEJRBGUw9pjlSJH9nkxtmxmr
Fdn80mlPm7Y8UZRQMR9+pAi+jbc0mezScK+7+kBN+Rq/WWFKjDMpvTTwMjY+gQQ9l4Why/c03DM+
Vu0AsuUE9pIZFzzrih+2hhLbdRmMm77vRO2J9sDxAZoC93mJnM0EpZZ0wI82N5m6xTon/7sbD2Df
KmdxmxBYecaMpffESAnCV0BMKpkQ4xTzPI5W3ram8PE9wIqAA02mntei/jzbCfLqiQUuSpITPqji
MmtSziMEEdmE6xM8clgyQV+DMdJgA36Ia5WNvs9ql3SI/PBGJ59SmCbVp72Fz13Jf+a2kg3T2fZQ
2SEm7n1/B1EQDmcegqqVm1B5EecA8zNfA3XMQLb7VM0Z00czd5YgdkS5ul7ItzCH7q0FwWySVutu
lvXLXpuqVzRtAWhNzDh5fKWw1bQDCvJWPyuKRbLLNdR5svp4PRZCb7P3/NBsyrZOsp0jIIo29w3r
vSd/nswVE/6v4US139yheMfDNtB+UbWbwkGhB3wf4g0mGEjGh/2frZNI4BwVZTumHkaWCpBA6arw
RIVsO23NL8sjRKi3/KT3megD5Yx4R6FA3VsUVWZdHBvMWbp/cIMgmFBysa2lLlZPcnAjay2L4Dms
wFAJ82zGG8X8qUdbE0o4Lh2haSAJafJYVbfHKLWNoHPWyefbVvHZpUxJsgcRcTSLJmklN4HIq1y0
htNH7oM+zi3tsgWLqI0VqAegeJl6VV6dOQKFJohAMI12xJpVBwh6+QS+cXVjGxD3aI5F5z6a0jTJ
wrFGLeBfgpvAw/HHmjJB1J4XxDqK2Gq5SZn1WTF1OVgjeDrotuCUACA7a2bHIZozd01FGKOvQ2Fj
cLRqnrdzAyNsCnDHqwuP20gEWv/Sjcfy35RI5OpR+umR/vzoNW890p1w1vO0xEueUJ8v5Mls85Y3
2vXBnwGe3ZxwIYxdWWsIA0KnnAkg43Z5Hdx807inyXPfH695Psu/obp9wSwCEfDah38LOVj5aou3
ltOumm/nO7HP/51D4XVyKhGjqTL2TSyXaZ+Xa7h7UE7YqcoqqTPcAJftSJHcBMB3do/cazmIKzQW
JJ3BZiDyLvqZJWMMYkodiwuhi68NijkCJ22/zhogt75DpLZYgquDj9aejHCMvqMBG8Sc9bWAuuL5
qp7fKDRiuk2bEiq7YDgTg19LEUlU12E0iKEkqcynSanrv/qiSlGS8Vx0UAu+3Ko93Wa2743jQblS
qljBYHm+28YW3PT5BQXQ6nP9bX+VEmtkdXvTJ6f/g9uDqeE4ojdBepkoYFXEmYenDP3ckc1jQG6F
ia8valHf2ksVn69BsQcsroOpkTva4e0eO3RXwfk375nYUO+n0KtznHdCMDCFl5JYlribIH4bCRAH
UWBVb5Iq7ZFTesnhsBtzT4BbVB37wJbPl5BXUqiCBsHZgaxRAF52yDYub8saWxL/usiV3rL0f2rM
nwi5H7Ql96bbsLYW/zZdX1ApQuPbUsX5u3Zu4MmrSZ9/+sZjZtMZnpyW4lXP3BAIOiRy390YPwhW
ad32tK+42TbWSyEwrJx++0MfSWQPDd0bsT7CTxrNuVrwPE5AdAdS6m8zXyDqTfb5zqDiWJNKMIzS
zl6EeN9a8o7pxMRe6Tq0h3sf6QZnZiS5iGkfIC2zMC5OfLdBVs/1ZSFnEXA8gv1NpVH1aAIjJcwG
j2CMZeccikaALmdZDUXKsQEBMPWyNZ+Hrs61RS5+1s+xjjNoZewGvf85SlaNM1i8CYrpR4Fn2lCL
99IuoHPT+cIrMU08YWM3JMwA/rPqtqs1lC3omvAUBQnmunyFglB7WSK4c9OUTSTeVBJANZ9Z2ofC
DSi/ZdIUnCwneYJl6ly3619qgXx5+RSHC7snWtSaASQekCDd/nIi8h1RBoFUY2FmL1bFDt3w6KVj
x4WVWnyFeJQmQQpHJ4p4cmtZ6Hyku/IY/ph2LI0gqBASvNQBVkA+SVnZRMkqvFDnHbTJ43qwVMNB
NfceEuy1IYJRelJhmpn2W432d4YVp2tltbWYPbwIiRuZXcBd1ri+D685KvI2In4P/cbIGUx7bCXj
mSCbwCxaR2Yn1rCPyf7y8j3NPkFE7/A6WlrrfdGDJa+DA9ZMM7khYIekN901XUyPoh4QgNEOnd2K
LBJV6CE+1k6urF/aFA2DhB2VOK/uy2jLQdnLhwcMH421kneisp9IZFP6vQjmWCIuku+v+1PPVWkA
1Fqi9zY78aiJVFsXEsydjONjR6A+YwhBVEAQ5na3bAVSd+M1e5bfYEoXQZ5dcoLqIOuBu1vjZ5gu
GElInyi3VXWYsZv+GdAz6M83cJOjoaEavnNcciEgZuVd+7wu8r7KcrsuNQCaXyjxxD1fIUwtLImo
rvX4wKMdjKISORGux2yfUYbU+SU/Ett8ux5AN8igCRy5QJjZ9iDKxCtUWYdR5dSM40UxheRi1sFV
w/8Cb1xS89ol1Ru0Lcjnoq5bmpLodLcXazXUHbK9hKcbyUU3rxpoQ6I8GGYWlMC6EzK5fgYJLCNY
Q5rJGmLPNHYD+j0dUv0ggy0beh/UenN5epnXQdBw9X7bdcfe5/850SV4oPVLzzih7sYK4BRemZLE
D2dUBqb987B+YArGeB5RL+84/V53w2XyHD3jFBxS77fof+AFNSZAP5dhxPGuaZsKHEABcGmd7lTH
GkrKEonJy+0lrtKglbVXc8Kso8Z6GZqdRlSk7DbKBhBAr8stVj27Y2boS85FoD0FwUMI+cj/JdI2
FY4CNhlaQXQFxA0pnmOwO3NI+D5dDEdtA4WGeKxJmowGf8u9BeWUkoQT2ugaWdUIJfdylo9dJhU6
m4FlchimRQYhYAEtpFe8N2Lp3/cOHtME4avrEEOk308o0EjfseJqh5EJ0dESpWoPKhF9+ueo8JwC
qlW3XufRpr2ULybkPJ/UBZZbYIkWMEUOVUitjkxu78KYkwaUJb1DVoP/5WpkChDlJ3+zaelRorMh
xrR0c+HhQrqHlusVvCpo8I240jPaFm6p2dKl7Ib01r/A+MUuET6OBmvUuRkpbSgFUx9ATSKp5qhk
WeiyNA7/p6DRvekXjGgJxxMLV/3gbLN6qkRCnXCKGZfUyspSn3vHSbmRQdz/c168X+gG9SsnuXww
HnwfVOJ1IjeqtovtAvSDc2ogyz9YIDYQuxLN7fnNWSuIFrgklzQ9PEh3UTIuvV52XoXlr/A48rH3
zL7DG6/grIcYqWVeeiOLfbzDiRrhV1k6vkJ/CCe/B3ASZWQO84Chh7zrqMk4tZRLTsaSqTd3sppY
faXQ+4TeYQ9r8tlr3u8LFBTsDAjKhQbNCCw3DKZqpW1ofp5gcphRfflYym17snsO//xICfF/xmi1
iWyWm525/evdJVVUqlaBju9ZQbhw4rBlpj1e09z2ovcAdGfGRP+n3I3MhE2l8onnlZSIVMlPcJRp
JPITeJ0nDNV6lSC6FG/l4RbDQZlby8wAiKcWyGkmmm7NfD1QeaDgtPtho1rOgehWincJ+kR+BRZR
ASBvLlp3Cl3HyMGwfh2m9lDHfMw7fBC6nPSEvXOlsatA+Nl/YVh3V2eky/JmhnG9RKj/4E9BHocs
Aw7ncsXCBq/26EZIg5Oq9/erPIN5VQscFbe4NPlsITp6UvTfoXRba04eZ/g9u5+m5urcYmolIkVt
pUAoXTjxhAZXEyrbOdXF1k/PWuMYUW3vgI2O2YpoF4lwEYnwVji4b7eUIq4XjILQ0urV/ig038aJ
vrmCcb7V5zw7ifmzE6LwkN8LLQ9XrllT1FfgmiKt+S0wHvoNt47jQsDkpnph64BXfGlyJ+jyLC2C
5QX0iu3ycMKwOlnvN5Jh2e8kBjuraUf70kGyIZ2ebKQcPlw+xCpsf7a1QgCmWEJtwO0sjDq7XT5h
NuWkkDHHw1F7DBxgrTLyHE7EB8KScswsehqgaRga8JqSmPAofDRTLKupWUU3prbYSWc6ujy8ffnL
i0oUnxWHU419v+b2pHfgPLR2vON1WMQ+gWg1KNEQcfXKTTV7x+mCiEeO37GJTw1JDwqFWBY/3rzs
P2pSV4OHeP9LsAz7rsLVCfENCgSWFJOVsrmiAH6qNpdg4cnCbYDby0qsGhKtGrPC0P+2tncPDrWl
qo8tgyx4yBBrQHPfJ7hYGIaxVJvZU1fQyK4vZPX52z+8mdAjqtmDZWbdHbuioO6LRbSCj7Ylw0vg
hbNpZToXKaIalNCr7w17UjoFJMAwhaVDoBwbpPYauChiFLQsNtUEEIGNORjO6W806Jc/66aG2HiM
54MIq3ET0chg7crN0M1Urpv/2tGfews/BBniUH2S2pz0nVRgA+PFnjNUa9HATD6vFzR/KALINC+m
EqUnkjeQmVjIIYgF4tEPvZC9O9vDwyDE2R7RMimXs5/bNZwQz2FqxFk9pDdNENhS5BkFeaplq62F
C2vZn1JxRViJDAi5S+hGV1ACd/A9qnY0dvfFek2w5N7P1Rohc+ddjeIWe3bWvM1I2+rx6UoaBz6R
nGLb7/jA2X1bAG2kabwRYg7KN62nkTYeEwad3WDFEdQRClCjy9lGtQO4Xs8iGRY6LQsUCrBENrQ4
FqqxVnWFjrzrYawpINxNiIr+T1bxDAXMCfKkSffzIn/GMeNw9+l8aZSa+Mw0Ofy7VmQYpuqcJNXb
Sm1/xcjFhlrVgM7EAOfudC8LQoXxpoZNbjEnKR7A+M9H/IVBXnHs0MdLQJGB90tvZT8WO1WO8gxM
nul9VaUIVeTlbjDTw9s27y8i86iNYySc8J0VC8tlPGZk5sm8jLP+NT9eA+MBwGtQ+HkN9y4dtJCj
cgqdH9b2xF8ynexYEVwZWtSU57MwFVl7dC3FrtMqrn6VK8b/tVUsj8aVMGPAdMUXEcjLiaPEiOD6
r8bLnxGlAA9XROo8RDvP+PRmXe5PgdvAprMc6C1AaRJ0n4CRxq8Ls+u8Vb9w44i/i0nlm3spanRi
xgMoye4bW7OhuGT7Pet0N+oGdOcxw2FGqxr2QcOMEOYJdIlSmb6TfDQS0PRRobCEIjx8Nuq169up
x9GEcQgi/Xx5k9PPKCN/jTs4c8MlT4FWKvbRjcfwAGlFf7P5gJpc+7eOfALWZqOP1QMhoavsB2/s
LfIptipWAWHWbFyNhM0KKKhLcB4rIwEZ4dLWGX0csAhg9b2IH8c+fahH69jk2hXYXoU3WWYZ1j9j
17R2XxcSFeg/DcVAb3rhsjkx49y+c9alc/5fec2wiSaKf91NczOZJseEki1w6hfX9517llIWEbn7
AvmRy7Pa18KTV0zHD/nb5QEuo+KfgBeRvJLyKvdgf5DxCuOUBb7MTM+VeIHmLQdvTqMmmZ3WZNxT
fw+l1gbfLYa6A71Wwpf1TB6MeOusQKFs9IJCzn8dLAMdR0V7AEfXl72HCxjrlza3xnbkucMZDHdV
4d7XtrlNAi/XuwjEIKVykGFQWi/oHeQhGqHHUvt2qbx51JVLml7ppJmsviFIWUrKNmvi66hfFLbd
FUFVY11H4B4ssyCZSiFaBbX5iADXjM+12EVePHyrLD5W0qKPV6qBD7x1bnEN8deFAZ1gc2cw1tdI
Sqg+oarUbsl5b1Ab2gSIu/+u0wGDQvNiX10NPcMVETnT12ecwBMUJVC4SbzPYHaEgaxRyiAtejY/
ExiZn9Y7kPvbIyz/K4wem2IE5o5fdmVRQ37K+KJpIIc0jaSBSQJNzAzSKhSXGwe4fvPDCzukdkMm
mTdyAB2CPTHMG8OtaXbsCcWTnW0+7QOmShZMbErVdLeF07gt8CeVRGYis7M9xuJVuiIX8ps9Ak2j
G0w4LfcP+IrXGzsIqhgrwYmvGxLFjDWrlmbcQDAZH5bBsDC822YZrSPiKAz09JewfDKB9xB/72PK
IggwPrvsEMwk3c9Dj50sTHd2uds4qtqnQ8xhm6lgOObqErco/QDQ+eTZ2eZDcKKHJ4F3aScNY8T0
E9ACabAvRRYGVzo1/7IQeRvq2DMCwIkKFPiPEwsb2zABYCDmALGJtZg2RrMvC/pgofCNeBDUz9e5
J5fgOwfhsKVao4P27NEQ1bSQpm+S7JbJOUiMuvVj1HuV6L6Z6peyr8SRRvCwwJHaRJw9SXGixK7z
qp7wBJeU+mL567G7ZCP1G5fdYXSlxwtUVKa7w+d+LYDPddSuiHQT4gnaK/XQL7/kKyRC5+AApt3u
u6t/bOQmcjTUVC9emmQrjayBBNmFN7oTr2y1c7+iMvd75WgUGbGTgIqESf+YA39X8aI32wbIKHrz
s9K/SCIKMlSsIIeKtIvo8AAWcK9/x6NogS7LKhuDHjZe+t1EpAhIyAh+VLUxUm3WSIJBvJyj2myQ
5kB0ObwXO4qzHV81c/dL/AEeNHsUHdZmvwC0zPPaL39+MFiAt3Sik+y/Kp+VlWw3mAeITiYHx1UX
NFW/YPnQaQ+Veq68hXsg4OI1+MpQ8z4N/cRzOYstQaa/Wk0arSJ5v0bHab1hFA5GU4qu6x4Sz8Kr
nadSN8/+LhbUCxVG00r/cj/pxquwJo3aVvqDFwQDCzkXbwX1+u7gZoWwOAiVnihT7AR9z5mLSLCo
APQ4NxMSR44dUqs/cvHmDCeuNNCNOqCjqc+J057VkyfFHkucz+pYPNO3uTFWuq3uNEb8dJCQITNL
akTuAcl7pvWBAVtTTLmSJi03ufbXJKo5N7irK3Rt6H0UK+o+0WWMbygHnumwjJ0Ys4eJd0v8RYZQ
rpeiE9CztYvCBBWMpFs9kYS4J7/lTJsEDQvu4NjwJpL5ArfT/E8jLus2I7UDbTy47JAVampUFm3x
qXa+aUIkMt5mWBNGYm2lHNW9Hy6kM8h0B0lhUWM/FIagqEFrQ19vBwKN8uGJHsesO8PU4jluWyxy
xjV8bDbwNBkrrevxZLmYX+d2zvhiu2XcNGRdFEgbAQZ+j871XtyT3pwl1HgpTkkhRIqblLLUj9bC
54ubKzV3y9pCP48AoARucy/QlJOZKTlqKXwHEa03NppVzUKdOr/H/k5BASEmhKJmWXJd8JLWQ7oG
FO3WUoeTx1l0Z5w47wbWnoRqeLHOfzseySAf4VLAT9MT/kRLTTGG0f8QUMLP4acL1UHm6qCxapsH
CbvU6imTCAVR0Ru35g8HrorEpEBOp1zHbiUk4Zga4O8YdHkNBYnLt2uM0UcQxV5yN0m0nWSpFOIR
ULO51UdQ7ws2ORKH3IZ9eDkAHXfNKaMgsD6zpMxTZLHMKtqTqTChCO4NMsLRjWUj8FdijO1V9ngR
2lOq8sdeKzGN6Luj1gwvQRq/yGPIjEm0HT5RSr+mRLZCTFWH9rnFVxdRrpiS9rebbG972dHrt3+S
VxlnngmX9/We4f/A4It1xErR+LpJVw2ZvhgC1lStf1lksZK11jFSs6QXmZM72rdGu/EZmxga/P2R
cD2ljyS7W/KJkwvfpA1UsYDRMF8X+XeNYst0bATcH7PpBPw9j3rBM66QbdOKyBVHTCjMGRA8tGwc
zCA/5XtGJUZj6yE4TI+IsEzKJVfawznGLIeub93ErJUcOZLC9SXLLCVW7+KRnhczqGRCzWVoXoNZ
f7EsRj3JY8giTFkmzU076hgG/9V/cI2ovuSj1VH7oKw3iWtvhqd788LAbc0qLjzv25uz0TnEPGLJ
bZtYfjou44t/Rcho5pcjw5wkzi4jqtPT3zCACtGl9IgkQRXT+mkV31BRaLf3NhoMozZYtJDeVXbQ
GUeeBmlCm0/ynNNUvi3W+sZ43zH1fAVUtpr/gJB64upVZKwshlomzbe2BfBuURo+5EWVq02kTBxQ
+XYAUm1cqtATI2yLNvqFyPr5sXDrOAA+y//z4OuRGpUyY0vaEZIPtSmZD3uh7OI6P0nuWecpIf5q
F9ln1pBWEKaSbb0jR6x5tRXMjpmwc2zIEuIhQxQxQ2F4CJHUjJcl/CB+97wzINOeeZARhvVU0Xq0
bQlCkoXAhFoP4D1EUQ8S5NSQ4+PGaZydNfQp3Uz/NOGDjF1mm1jOmZpkGSDdCUk1UQXYpbwf3gKX
jTtGtaiIr6bhWBB3RqTyn2sSBw6qhSZX9LlJH4PWhoOFDL5LTrK+aFmIvz5WiVRao42wZ/6vEoOK
sC0YPTFn201/42ehSyRevf2Mc6wiNivifKDNff4B1BGMIbFzE/M4xvfhjhJZgP/kikZpimobbMiW
d7kQbDcHnJgsg6mSE3dAf5HlxZmGTn2RbS3h2CRbSSIBdm0IHBskofQWdZBftd1hlsIcrOPRoDTg
/94MxTWFy/FOC31GsVVJ01D2pO0+gtGEYY1bQTFcsf7s7Ib5zpAvFTtIabqu3ONX51t+rBEnh4qh
YQxZAInOXAFH+uUZZDBQXN8ocks2C7bfovs7vlRtMKkFL89ay7ognf1k0eXkrpL+EvUSAuaeONda
7NVa4oohldLgAzHWaulyg4jxVRnKKq7jEenbiE2+AzRcuR3rQlHhJqwVj4otg7GlhKZUQoJZB+Xq
owHGe5LZ4rrpA4391QlQIz8xPNBK5C45qiFCNjMObW956/bYLyu/wPMx+F8RKcs/cS5TfumJ2p1m
GPHiFyqX8HLRKok9DfWc2NXG91S7p3H7iIRf0XpXXof09Hmwj1ahvpuWNWNM+P91otozLtO7OPZY
q6/zt4bz6BwTmQ49z8lKyGfaW78A+qVTDSFY+/tYrDOD7rakIbwU54k0kB0G96QQhxVduMYgclyT
23EXL2TvUSBB4HkbVa4TEcfEZrmUts7qiLoKxD+PRptpoASc5Y5hGb/p3f0pcbo03qNbRnq1hU+6
mWXcfy/2xC3UcChHWQAkzyfS7qkI+TUbovCpY14n6RsIm0ZIC4gftmSfELRx9qbesUXMIAlPsRT2
mMsAa67U9oel/1VDMyQuCP46K+hbwg4ZOxd4NN2Pj3CoP03wrVC1O5v3CktIHjOlxW+rF86ArW/E
pxRkwfpEtQUqIbNzKxViyInOuJYXdKTL6K4m8e/6WD9AY15fbcaC41w3naE+RjiTpL+YNVfyKDr2
CGePvx8uJWmLEh20rpM/ixtkU6RneQW3BDIZwgNg9RvGznQ7KtB5P+3Lnxwzl+LeuA5mMs6u1U5x
EnIW+dh7/8x3FjFiPZGOzCJgGfWHGrSYMhJPKVqrH6U1Ls1NCXCryg1SFC5FPWDkj5me9YUQBUSO
alzw/tNlG0btK3yuWBDsjnJo8cz8qZODr2RRFQOqqTw3i1m0PwJFKy48SCy4BPUrtNC20uHE4aAI
p8NCQq6Ajc1aMBEq43QX05LnpkDDdAIqse7gH/R3c4OmDF7uEZJtP3ZGS0OO62gcZp7xaHKPDH5D
cQtwzpczfIsK4KQ+fKozBuWTo/JiRbL0ODugtABnD5XoUrDeiH1q20j22J9vL7oA8eK8YmgJvnE9
dUghPbMJ/xp05h1a4+qvy1yssz6uwzwgN0vF8mQ24QvsMzQY2H+DlAgPfU4Li46xNeIDDlW01GEx
c9wZFTHHJqkMVkSZVj2NelOKdTsef++eI6SF3Qn5CPmTxl6KDLcwVw4DMbRmW44AL5ncqt8jcMsT
7LE+Ddw1emef/MqIk1qKAsKpQhQekQ8BozWp7B0Iy2WukECBE5hS01vou+vRs0n0Y03QdT2RCidF
1Q5CoS35ZORVmWAK7op/PNOqTH8U2rBexNmmL9pFQEX834ZNUGBqvkGQC50k8MEVeKaTRItBvsNK
jA5NFCZyqvS0itqNPameVFv4X4sFxOZIIXwhxhu3OsIVhmqWWSs02wqGdkOe43Rzz5NcYQKVej/X
+qcQsf3/K6CBWQLQk7Ka6awoZPfU3yTJ0SXaJXELGhiH3oQCTcaWwW2ZxPvwQDbpw5JkfF40jLvV
x4eUBA3O2Um2AkO2f9RBh3Byl75UBjpJ7mKFDWjQYZWN68cH2/95TUmLwig894eugRkCrORNPeIi
Gqths5KTWZ4ZsKMm/8383Bxl4N4zlxg13FG5gtlGpxwJy3e5QRMtoBhqKo/ruseDYBvYKOXscwn9
puzB3E3SA32rRShE8CJqbeXV/0OUzNIZIpzMCYzNGOJp53s5fRnu+p1krVRgbqhMlety3Ob26q6G
M/gNbb0cOWrwoMGlCfkBJ7QS0t5e+pEUf/VjancUSS4d1bUWdGuAhcK06n7fFL+qqzusDTNNpI5k
QtqUhg/yhqKxoHhBoq54JeiiANg6RgYCcUv5qI1LmSPOjANhzTNsKxYamBtoTzT7bC9b09g6xKQM
Tudb/fY0vr07S2dggnKplRf/+FLK7QHrKLh6lQteIY+RAjH+1vZf9oWZsHk01ay7tJm1Mc8aygib
7b9Eh0nJzh27u3KTjTUbOJXk0hes1hdlEIBrqO/08m7bSKkV/V8aUjBy5/8Cpb9mBFBbUzwdk4bJ
vwLRPl+bEKtMrKdYfgtWXl/Xh153YZqMyOgXoTHv61ah7etowmufUXPRSjPgvGwlOWGeGZM89vyt
CNw5vcnHL1xTjOiiIeCk8V7P9Vo79VVC6L0FBM1SVkyanXv1lkeTfMCAVNbtc7Rauud98hJLhtAO
2gmjo+fYQcnPmOYHnOzYMeX3cHscKsE209RqUqVK1xJ0p1omXjyGmgbuqUS2+JZ6eJj13ivoB49K
Jon4cA39c2Ec/ZqObIqf2x0kKd5KrSIM/ZuD3PYDJh7qus/lruvnGxI8SM0KikZ0FKYAArD74XTN
KM+JqEb6JMTVdt9Bmo8NIlrlXi3hqIxGPUCE5WMbSLdgtBzela4voDJydgeb1D6SDYEBYZQXRsF3
mwYx8dpn6bPdDnyFWghYh+PWDrrazH4VX4Qzben/songrmMgI2di/SJcVpZNhrET3DiCiR6CgBox
YEyBw7HfRikh3T3qoC793ciUpjUmlplKT5lawalLrO3imKE8hxLzM01PxlHcYJJh/b8rmD1JA2Gj
SvelBEY08u8OOd6vkFrqxgydZjQA8qo+1q7rm/1EN8bXh8brFJdHBL1iv/lhB9369HHAdU3Jg9Mt
JEv54OJLrknAx4fov3Q/EaxCD40hAr54HzaPvHQrdaq/Tdn410hI8l2k0/JKUjN8icoOT62oPn1j
jQNH6K69tswggkmiuDdM4IGw3ToznDlEnK7rweb0zE/c1dhWe5e3kQ2lSMfnRUIR+CsiO3Nq2p7V
K9lfbfYZ/5c29MHB8LQzYTgiRR1ndPoUgV8gPPtLTUEN8OgfJ+EzAQJbId4Ri1NqigxyitY91tnJ
HUAqKEzS+cslhxaNLw3IMVwbReVpNocnySJrNSb2jD94/UhhKWvN9H8SNFB8e8JbQ3flqgjIXLHa
ig11k+AkDyie+yeUIAQbqyBWFUzFyLFkyJqtVK+UubH/JCl80PwQLe7J8+ZdzBm2vMdmWznx3q/N
NCiOxtEWLH/+zYfnPbAXe5UBL+v2pwtvoXYxOzpGFY0sEwf+Tctaigy0K+UyTdeYKZ072oU4LU5L
1l83jBbZgqAa/LQQce/33Pu4x2O4vuoJI/JeYKbPcIiVM9hQ5Gzh/FqTUEjXx7D88Mb69mdNzKtR
3+X2T4oi0lKyIzx1Uw+iPJvWWtq/imjW3v/lgDnQaiJ2OBAq17ulMJDGEwgERV/Ulo47GClfM9yX
/Y16n4BYnK2s8HfSevleJAU+BFF/QFsACge8YprYZm2qofY/JLv+fWKO2bKV6qzfybeerxiraum8
dhwrmkmMgrbEIWsCxsMP4Xgm6QDeX4o7P/Vjhsrvv0k6i9mGc7mWglAzmsuHR2TaOdNNP/c3quBu
eCpvKIlNhAiV2kv0uVPxbAWZh4rEMv1TEOckuSP++0wec/qm7nExwiihgNOItLe94PBqXBiE8oto
cFQ2Nm5DdVSFt4vVK4WwmVkBOcbqy65qQzBDgfrTvZihDt51oWyMx+lIm3roI7yKyhUhGZObEccw
o5268ykchwCjJVSiFe63j/zNVQvfGK9yGthEL1C6JGcwOfPjnB7JOAxSE1a0yHIIadHFGBXxfUci
s1dUqNLZmgecXEiNOABjai4ij6r4Xq7F2UxF+uJtK19iGPiyoHcGyoO3oHzdt+imip0SJzplT9gR
GDMaG/URf/uUrH0/EUgN2HD+wLlqIaGfTLptWkfgNlJP6Z0kxQzsLwOrlxddlVl3w+hpoZlCCUZl
FlWUP7nARUq+eqmfKxwrRnVi30dxM57iVsqKCgh0tMQTUDKfN2Pad0xvEGaBjI7jLUCxdGXKbxVz
sfzFHzeleEND9UQI2RLOZnu4qrIJWTQUHB0Mf9cioT5zLLwp8Hc2re6/dPUc4llZ1ZOXlFTf/ZrR
JxPkBwoYfdKePOqOUwqp+32sKwEMiK72y0KRa4h2yPuYuHvI2ydsPLU15rYW+83QlrE0eT32M6Y1
8aOFl+Dx1rMFvlfN0uw7Qsj/UFjlmiGLI1AyL3gUAkazC1kZhUFYR7I+Jp59E17YQqpU8GmWf2y2
X+SmnakFbmJmyzocgGV/kzDnhDjxLh/kWI9Ko8sIVCL93ghhMJsFcuZJl/XT578Y3EVAQjfwC65h
qzWDvbIrF4IkZsLuGmrANeKBnmAdcWtBc44GuSNIwGpqLLUHfuHI+qIu+eKXLmkm7LPnQRhR4/tL
EL4YncCcBi9udBq1UZwtBkIwE32jAQ5BxB4zOUckuR7aoR7LMwZQ+vkxLc/ZapdIzp3GqY669I4l
HJMXYJCFS9C1MgieRjSh62MLGmv1bFmHYDYwqBspZXsYP9j/4PdkAiTEe2NA92WiLbs+BOV+oijM
E5gPoPTORy+7e17QNpXD8nHOey3I9uaIkXDYltg63hYo0dX+gA9XmioqSbNp3RUJaiDlpmaFWVq5
U6aJjJFvTFUaeAJsqrc/WKrQch17ReGwTg8Io8ZF4oYRGXl6e45t9TmjE0qwpqwAfEzDZHyQcE4N
VxCjW+pFP/PiKnFVKieo9i3hZamhGiNYZdiBDZ+ZXLwTtjYVWMhkKgBgBhvdTmKP+hWtdyzmG03I
1fyRumDHj4kdMHLgYrbQaEF0jymIfmae7thgYLSSwijDOJGYAP6uU3+AB7tXsxmLP1CJZpO5R7uA
jdGO/83qIPpRUDB/bvnmE5PDtZfO8+vLlj5edpIaNzGCHS7dy3srYJwk9WsfbYbnWR0kx2iL17hd
QkLwOT//8JZbJqdIMrr+OZkef3O+ooYLpFgJWTFeyxkes/n73p0oYOQtLGfth1aefzLlONwZV+sX
Zs9tthoEHimB6qFOW4cFaRH3xPRyzCME/nfo27fhniKjQ3mfeRi1lvS00efaDBjc/ysjuwrXRyt5
DMNSbF8oMn+Sn0c99cBjy4BoU2qY7VD0uU+phhiObCvlriIFm0jUmPqAHBAYxoLseloguluI46fd
P2LKTQI7qSvvLHCA7KDwANe3btbsuZGoS1USH8d7onHMsNuZTN+JegxlBAUfeVWfT/+n5scXYLhC
zcXDpt7yeFG/cTLsgdV3QhAANwuACkXzNgBCO8oAc20QPWopJJSUGjD/hPXWyNENZY3SjmJ6T0LC
49uphuUZm8BZoHY/3Fc3gRoRlqkfEdNnqrd0qmpRvBNzi4V/qYFGMZDo8ouHtLmHz6Q650WSyRzU
7dpx4s7akM0XIl1CBmWNom4apY7PjG/BD0WxOaib2+cRId9roUd7spUy+LiXCDjjs3s537eSOi3l
BNNxpFifbKO4LEiUiKjJMd8vj6p/AZh4beI0EGS6yIEUjSe0SbwHu8nXyBdayJw/V/Z7C9gF2pRX
qXg8p+kz2HSZZf9j/pifbk3OnUDvUH1A1PLyNas9fF07gtrseP9+uxJx8AXRSKW50iRLRyrCGpvS
sIWDnu866yYq6FV1HkUXLw4v42YP2DBDHn3E88UYKigirFR73zqNuy79LDm6jyqe4OSX/pJs9q6s
WhFDCzqfBUG6IBw2twaMNvFEHM32gvmdr4alfA4TdhtdoRpDYmHjYyvzwBkrEHjBf3yLqGXxBELe
ns7ivRiQG6QSLzMiq2OtF6Kxr2eq0NWUpjSyFiH8xVD16dMuXUTFaiUouZD/wgVexOsn6ONvDH5N
RKJ0tM9H71PxUPCmq0jsSlvSBQ2gjyrHWkWhyLm3VyNTinayS+k2RxzQ9iGdH4IhgQiXx1SiV6PV
cssTHcvweX9dPkFam6Y6faVR6dfGTmyUI/UZbrIEnXL2tAZt0Ro/HIsMCfGoUZG1ywYdFYOW5RfU
fWvy2Cq1/5HiFSQIFT4o9blIKRksF3h63faOOelAKYZLDWNuBHiHp0qVUXp1eqcpMnTYHbijTCC1
qo1UF5Fvj3SVrOKtNdx+AQq8hKUnN0TIRatSAy3JOvckCUTO2n16iqeFXEIYNXu3xK3mNnSBF8AQ
PkMqryNl0qadH3obTOiNXnUcAZzwe/NymiIktOVYBukACwRP/lXhdBNZT/4sJlTThfnk1pGMX+BC
nDh5rrS//BL/5r/Epcmt5j058/vnHcA7y22kWe109+rCEDLgEPcZaO8I8FWtvtQ67w9RJLwhB1UR
xUKI/xzmSnqeFJtR0vEtKjFWDCyInfmH9oObzMDgfARVEA3plxkUldVOV4zZphsCZ495yn8mzZJe
xqTv+aly68kt9aoGhedDa22VPkKiS3shy8DO7KVtO0r/o8+04P3hPVN71GAEnXdaFshmrS1CZIMm
yRYJQaLBxjDim5WUkVXa5ktv0+TdMw7ey1BXVSdN3G8i5FYKyuvb63NGtPEtR3tDfTi3k5RfroaC
C3OAf6TELtXRHbNhB6kunpg11OlX1m/Tm9kRdO2AaaZgUO8wGgsX/NiSGPR4N6jkXvI2QpVaQzRg
5m4yRxrBXH1FlTBXv3hmf0rpQ3wcYNjUyDd5kFkETPKFx0HXl9vnZk1rzlLw1VgIR7irI0DQ3HTp
aS9CyPGpQq9LMiHZKDyVCXvC5FPMhB+AAr8kRwndj2eoioaKKkdV84eTVwUf/QB3pSCyZvkSTGpV
ZxYHybEgBeYsBqMISeHd+pf25C3B1Nq8Vhms8cpCN7nCa5rUGUgfOIZhji/ocPCDH26ZBC5JWn8X
myk0MQwj7uHh5hbYcsM3i2e45O6WkJXNxU/DqLeU+Mrkqk2O1/+a/4Egoh0Y6u3QCH/IzywepXkV
wj3N2DQnyMy+hAF/YtSIVoAp0X5lTklezr1pZJgn7O/iA6+9oH/VE21EeKCeBCoOAauqtyrp5cy7
9zYNJDBHn8qCoPQnhC+R9xWWgr22oMvpNeTuDe9Yd05wpeTnGGgEbvTKNOMvi/VyDK8tqexgn9Ja
ht+z5XcZpNRBscNV1DAVLMMkyQfl9s0PdfeFn+TGWC2HaHGUoOGSjH6AUu0Q9ZuQS/9bjpnSefJQ
YcN1Fs8J6zJVebGuxbYS6F2L6jp0cyuNgbAo79tl5+G7Id8wySo2BFmJ4hvx8pN+I2pdyPoH4kl8
6tgwYAc70FYbok+66E2Ck94OS9/yXynvSJL1RvbRjpUPUoNd98YwKhJEfZ7JflKv1wHgIvUikYq7
CwtuKL+szmbTLjpiTbA5E9yQjNHIZFQ0EBz4R0AHPLo2OsbmI0IBJXQEvHXM0A9VTwiC6YsUd7sE
nr3k7SYrzRSGgFmyKPa4JpjWnXRvmhTHLHsoOV6hjrp3FUBgqOCjouRazuZsbmGEKZqlitRl8mtd
1vG6Fheakll9Ox1TQjPvuIsJtLN9nBRMW5DozOd0Sz7DVq/tCyxXh+Tnxy2p8jomHm3T1bLx9qwA
UHqHTs8C6EnZnuDQKZ9wGe0d7AV4tInk1sTL28+87aNF0yCTxebxln5wZwLnnBzcsWsOIlEpNbqg
/H0Nw1H/CUqLoDQap+LubuRKwNcEk9SDSvAtmk1cGhdE7/dl0DvGY0HMLOP9i1tb7t22OA/ycPf/
DyEPhC485FAJpPQwiKOet/jNAc6ccPhc7xxaaKFPcBVjwP77jnxYOAb/7Z9IjrPu6nJ8O99nwAkR
sSqfaRqWdsqhwb8IGVDAu9BFCqaTOn2a8IBvmMsOT1CRh8wQJPaDbewCLEjSGf5vrzQ8tLBiFYcl
NB40nXT/FkGJsNKTSMoc6jB9npIMsXpRAunr+bFQAccxS4FcysF7bW+bGlubDQZJJy3+VgIwgQpp
rMZOJazFE/ogRgY/9Ky/V/c7GFfKELufCHmQDnmUPBYKaE1wmxmqUkfFn9yNnPDfQwXaCw+su1/G
pPKoivMulTfLTncpkUbjyYM/+I8YtOW/iHN3HRbkTf04p587C0n00/bcaPotkX0gt0RqTVfZcKMY
WFLpL/lBnwsfmzhq+7svPRRjLCPmQxAbqBiHp+hoP7j/1aAfySRwqsd9wc7LlOHqgAk5UInc081R
JtJPRnGGwb3auxVZFWlJ6TYM0VPUsQxgrfW5YTbNezVK5SbDVl3nnFP6YhZR2oLdtdeMxs4coVwQ
HDpvjyCzAVV2qssVHhJaj0XUD18PKo2nfYXB8J6GAA3hZtsxks5Uf3dqrD7+FLVLUdq2lbLFoFo4
qdwgD4XWyGCqiRDSGxxhn/Nq3u6oXAqyWs6J4Lbikc7VQ9i8y1Gebj0ki3aImncDseL3C8O7z0OX
5aM+Gip/AzXwKu45801K8dR0pBPz3xu4kzRvlNK/9nyx2O4FP+a8TnZDHXwi+le3PxKcuy+Y43h6
sWgnUrhLf2axGs4Sxnh5ty02XrqWyig6gbRE8tTU22a2xIK2L4HGBcK2ubQAKetuIf5ndvtt93Z/
MAFgl3xTlbrwsbr0VAY7BzN35s3jeyq+JpcPfJnEopESfgjaGnRyBSk3miuUUdu3NwUo7OKWkNA1
BTjY6aLvXCDR7MvK9GwZW0hjX9+HEZV0PloTVOUYXJl2qQcL5dyc8uYljRUNnuP+/IciurJMedBq
AZ0Bnr9DRHfhmfh1u40fmSzJOR90vtfoKheFbfMe+kABiveNPh0TIWSDJz8P04EqzMGJwTuvdwGD
sPXq1H0u6/y1HVLQvvrnIdtnHcFeuBz5PSYlRSdUtcnGOLjdRc/p0LS/px2lDWkiy5NdLVcpOTxy
5DW9NECjB+a+VS3fJhk64EZ9Ph4LuO16JH5UdPBOkGnErUFwxM1tcAy3MHC4Y9UBqVbCCnJR+MQh
zrFXp56RyL31qWhtvaW3XkNuGQTQcFf75o3WCfqgi0e49uL8kzvQuB2oBNu/ZiPtlAj64t/0o+pS
YASJhD2pCCXEn1VTg7tmjCewDj7ayOfJ4B0I0aEEsUeLSMI4nGOf54JAFQUcihOozpli0h7cAYz0
pr/xrdoh3pmNqFgwYeBU3aqhBTcTrHd4s4qyHAY+9fYqD1FvK3ZYC1o/7DRsdz/6YACzK6gZKKai
zgHJnoqW6c73djwVBX8j7RShrUhyUJioSuS7ycEaPt03blPAAwTtkkEW7P9oAW/wYgO+gKJEXvY7
OIl/StkbMAolmJF28pe0oWzsvbEQ9pAzKhPPjjTaRhU9tdJ5cQlFd0B9hlYeci5hG5ytF09CJU3B
VHOgrbKClxzQ/3Kx9UIDslb45bAszrCzK5awSP+yGPDADC+Ukfkqw51ubAR2tYVziqjB0vqGZXBY
EPCXood7smUcGQBsG4/HLLhPSyA90gW1g7VtAGAAMgru/NemRB37AahbWiD5NAugnmzOEOBPY7+m
losE3PbXoxmK5J1cRBNkkysg9/FhaoVf5sEGH6VyqBie7aypflr3J79GKBpG5NBTwmJ91RAVx/uW
qvTjkxNv/ZBP6iPknkLq2WgXcgbHihGAqKPleSSb3NRcEdATKLsDCx6hozKJx8mXUKNDMsL/Upbx
s24LI/qhZdcavTR/Cxpn8eYnbYfR5K9a+8m9aPIFLjh/sIsMb3hzM+AQlQlIykE36ZDmPpzBeGFS
T/nFfeQQa2ceoWhjmsI84JQEJGnkWryOg0Ce2GQHkza7YVp2cvJOSjssxztksuIKrtJXnDp7I02e
2FopF5AOksYMRZC5sIZ6+gHTrsNs+f3X64w+Bb6lkioeEA6rXy6DCAikQKU5zST79+xfVnmqgjne
6qiiRQsxmevBLXVXc+XhdjiqejW/vb0ijadaQWn6gAPoJhVD033KWF8Y53Q1Gkm/RhOFMvAclZIP
QKCTqR3K1kwMXZFoeAn9XIla4obIQ1qtlH0YQ5B6GK4CaJa5DkRSN87wvV7D5io4HZZh9ajx7DDr
v9XeMiMDL8hpROzjmX+yNiIhRYd42xz8g1wDmGnlTp813HP5QsZwzjsRGocNIcsV/d8PcZ7eD4q9
DfWg+46Qlivz1SbiQ/JuWkX5Rb1jasgmDIGjZm+g8gGidAO5Au9/a1nz/ABpAUKuKywC4yodFAQi
rqs6tBl4oEOCjoXabHg01nIq+qQwaRgUVArSjWBqSEahRZsysB5J6yf4eJy1DNCt79XqlQpmHZ/l
1QjtJUl17LS8O5kx03qVMbkCJ+cs/O4ijkwtZBXq+3NN1WDNWWstUW9bjLHhiP9x7h91/XRizFo7
O/GkcMVkdnemkEpvBKA7Qm5UeKUbMoOjVmy7cx8U+q/7s/8EDMeEM44Yq06vo7ZzYPD92SYkmfkF
ee3s+VQOQM4WxtVDErJBep96esiHm70VutGZNmHCZCo0RPBsZ3/A+ZauBYnxEsJnYtGmI83wlpxV
6ili3UhSx4WD3soihCWnmFoONUATe//p/mBWUeyF203081crxqfaMHgafPpULOpsCvB87OfTwlE0
Cbwo40U9hNRx8qiH7ooAzdtJDVEBHkMDuaY0jmLNl2wTRYCcT3mHQNBG0pCc1qMeok0o6XNsfxqa
RO/Cqv7HREL5N7Vr4oNLWc/M2vzj5EKdogmO3uc5CqSA4hytljij2Nn+N8WbBQVgZQH+tPM0/pmk
P76hoMDgHrRITXT92148rQGnw2m/qbnhmj1Ch5oS2x1WU8cd5JunHluvMxF3/TFKhJT+dRXl7vUO
xkPbPgi+bPHcSgMP7Bjv1CX69dOb/SH8Uz9EtTcvQkPdLyNJOXtU4biYSamwwhlj8psxqV03a5D2
6CyY6i8B6nRYs4F/uqkyrVQ1pmzXO+d2wk5hsJerST/UO+82D9O8Ejxwdfy9ZPZzanhvMBb00Mp8
N6n86fl2Qnz1+uhqPovodHRKQfNh9vv0wK6+ZHieSmwvtVcxDAMwCQMFrKpiMgqL+g4OC412XzEd
QWa1zn9ERdF2sOQ66vRBawnO6yclXdl9IO+HYi7sIa13/ztat+lPRY6QIqZo95zCBf1ULSL7Q3aa
mT11F/Fwp9jYaL5OqzcSod7xuXtFSJqGh35GN4dZJBHFoZ8FTZZPVf4HtPY4u/U3/ehIpsCUg58I
TNXKOxkvyQ4BYf/bZh5prtwt9QThFeHHNcAqrUZxULmm7v25bjhvwBHNYNqdhukuh3gmQRxp7aOL
g1dgpqxAMEpF14p1TTsGAj5jweE7bhZR1Lv3tyox6OkLwilPslO8FpDX0DW4KPvizMw+no01NjXP
jU+lFbpIhEGiSmiAruI8bSRxyVbYQ8nw5PptoOMaIe9OmtbMd1aZR1LOQLQIfPvBftJB+jcs36aH
dvWroZvZh5g0GH0kCr1ZuPvZRWdVE1c91szAn5wYXMKiOd6pHEb7dRBW7cEMPWPULDNDXmKmg2JK
loYp2zNF9/ecJ4aFb+AGeJldoKA9ZqHDeMlVg4/5AlbziVk4eFRIL45a4M2HgjoOArV6955kuuNT
AMEb+qBy488uZsCy0RbzKaJD/Z6zyz3asi92qJrDRurGcMAqK5gA2vOm6HpZL8nU1SmRUcNwzKVR
9IH76h0FXDlBFhy/1BJkyTzAvsX3CdVd/K60nUCmqFDHjDJSnk1IuhrvGXekgqlaUhMh/T/m4pjZ
4rcuouW5omL1nEOXXAXH1Znah1C2HqYX2Yj8oz/eEtULulqafLVnCrlTrJJ4RhpH2jhqv0OuE1sV
blZIE7eOojvlX238wyLqYPeJdrNPm4aDWygsCxg7pbbejPGD9c5ZgpNBUsYp8xWlR+zOOL+DojPn
IReSBJ2fQ4uiDObxj5yY6dwmWm7QgIgZyG8ykW6YcaHCZaZjFFFNCraAsquJXJ9VQC1GQKXbzQ1E
TmpzQ9jSIC7GjNTWOILDEEcu+dfjCaKaZG1O/qY6lOiU9JQzSiHjwuoqmMPXqmgHBx/y0e7hTpg+
3tyArZwINYnrlsVMoyJTJ739YXH0CE1Pc1euuCzvDHPh/YLfPZwaFicgK0MfwYZyo3nJ2fxghDjO
SzIy/B578Us41v3Jkg5XMSC1V3NeeZcj6nhO/MN/98K3mIWjnIFZNF2w3lak1z7lHR6kAZIduVVB
WxX1vFrXx+8DHDlPqUXZprHfhP35pI7utYpu6H4i3ydQZtVnagujNGVSbphFraWvRdeQauQqLuvj
0A2OKzNCEBhWYpsZHDxd3Ln7mTDRkALiX/lnq1iQ8WcFP02EO17ccp+0oeFhB3jv+nd6FD4PRyrx
JdI122wH4NFv6ZUqPKM44kgTJgOvmzBXTcOhBxR/8SIv1lYYex3xFE0qkkjh3R2IpYYa+nSItBqH
kvYigwTEo9sIEDKMsN/gu4vW78Q0ulsbrzgINhJY/D61pHVWoa7NNP/yeJOKTdO2nYcWqytZyY88
9TwT8gxLD8FX6bkfdyQJAu44am5l5TelKWaunzpR7nVgT8SnBzhBcP662NYOC3PyVvOgon0g4azU
jIBe/8PoNFb2vGfA4vesfKVu8HBNl8r5OuYaJPrf+HR1pv1eTXSIfDD8E+2NTtwPH4+7iuhHL//6
ILTykNru402h7D9R9XbMZOMGIAA2ro9ziN6BR1A1DrqraFAVU/KQd+AjoK6Nw1+ySWxX8/mmrvao
vThRvrHk4eLSTgcpwnN+qLutzo+scClOl3tdr1r7fsSPu92NC0kpDVqSs/oqHFR7RY5QbJgejuA0
Kiy05Ra+j762SsxK55P7ayluwO24ljriMQz4Hd7T8cBjzMbQFZxb0bd1A0RpdYm45YXce+iF0k6R
hhbYdGrSeBdgQ7yM5UODrouq2ds0CbAP9/2eil0/D80O0LOWUuXTVNnM/eTo+WSG51uQKT3opF37
O7aPE+iI8igiHjApF1gXh7d8Ag4HPuRIwAg+i3utqn/7emS4Cd8bX5g+1zvHV+a4mQEgcXP6li4E
nq5pYFvYjaUdquMe6gUvnVVeqpmMwyoWq31EgkgPX1YO5HFLEF0sWSM1Iw5C62a1wSJuWXQg5Hey
5vYfg8y/Vcw7NKcY4MoYzxcxHr9CXpg0ylGHg1OoaMdi6KKQzJGN1zJ8lSClemmwMfewnq0ozmg4
2RhXlNfNohQTa0ZARCTBJjId/7tJ1FVXdmDMOVABcCfjddatiCmoUcuxsGLG5tWBroFV0medvDZM
EGF3ekyqqgOokY3nwLCJ2mirG4yCQSwma/yKk7ArThXgQs2v6i+3l9zfOyKC3M1r9Chv5BYYfDXY
cQC6jksLa/s+pcj+ILx1EHLO3va3s5Fs754NKQm581XTCuaRXMtklYyU3r4rrs1NsFe748nDW0SY
cpM+g3dzEVPMsUw1ZUYukpwgjhz+zJT5e0lPr/1Bt6Hu8Y3BUXmvpYOiF5rd91P7W4vNJwc2aFen
vUkxoJOrSMDcBU5f777RL8pFf2DvfaScmrHwu9lhUFtaJEynQV2MAt3+/Y7UcAPB5y3QqIkOz8xv
RRNVkeellfAzMxAxINIad/DO3QZqXlnUZ3yi9trpUWfTQ78G5XRpjwUwrsX7ul27kjT7XZgWoJMZ
kBiHvpoTdfIrsp/rzvCOuzhtyT3TedgC8A8QKDYey+U47yrftwspe/uM1QpILQVtR7almCwFkQ6J
elQjcpC4oOwWJ+TCrVDhhJs3YXCRSWH7TD37eRAEnj01uzLNOifQiJ3yTkic+rEVGJW1PpRv9q7J
b8hDNMPzKQ4BK1kusvqPlWGYgzPN9JVV0tBZNIxx/xkEP2URZ7OxVrqlFInYmbpeHZdvTDtLdR/G
VvtlbhTjgXgKJML4V4QySvMCT2im5ehghb2awAVMmRPQAsZ0NAuAjv/fxHiTUZQOKbPMQtTP8WFc
1uvQ8wX4w9VZCgmYd2AifSjNfLbJjzP9bXFniU0TA6e+byVofAag9ksfj3OyeleyryTKmJ0jSczU
d8ZTsDow9Izc+SNzY9ZiLE9qkHSMztz1h5WLGw5pkweNw83ksvcd/+kgXSEAVIFbMOj0BRYF+WzO
sgMVf3uJP1VFWEaXBloSGV/UonPxANaQFoxFqG796LhSXvFYCwky+p35g9SLbAqAckR2+JjmFJ1V
INuClnHt/4caWZg7+ik+s4M2zZsfoOG9vOE068jk2a7EUFM/TtMDkYpiJ+Py38lfhXJaFuHIcrQK
Ltj8tmFGLOQQBArg5f+8qUT8vDjBFAgaDp7S27oAnY9vZw/cDrZlhCvZ+H9+rMbRawYVr94T2CrY
eXu3ojl/jrWSbAgdmt9ufHHVJYnDRGn7c9F1ppdyjVm/x1aBqWDQJaKnNpRRqSXTt/TIn6dzdle7
KwKbI52BkIeKtkU2FrcphPFVR/Qp+GSpVKqpOdHeTuhpzg6qrwSSmCTSpxSYJfdlhJqlEGqej/ZQ
87lF6arFjOqhd2XvA2Oryhmvr5HvI15VYbHHqlRzyw9rRwvkgiSHJLXV0qLsznJ6U3f5ln+F2Z5y
XsBZYJWU5NN1KT+FI8IYmCUln+NfGn46VZYFgbREFdflowI76pWvQPlGNOWyDAmQ8iwEsy5ZKhBe
OV/A7RDWPN33Q+j9f8YQ8+NskcYpToiy6db5aWwtwSvKEhp+LM1D2xTyb+6zK9PvXbjolWj4ZgRe
Os2m8PgDNps38h8JuoGZYuyF4wwM0dKhamCtYGR2d6ZjEvGNUwZRlf1vToiDU+1ADHKz4WNFaZkv
YbI5YWjHWGIjvV2oZ1lZRFxpzGJn3Ti9exJfT9rGIadquYWGiS7iF2TU8F8XItfwnLmqN10RVf3x
FzSJzFKIoDNQxVx3zUAbAVFSAGLDtwHfj7Nclbd7jMrMMUVn7LLccpDn+e9K0s1jH3ZJQjerjijO
eWWP5etdVTboiIhw5htxQwthoFh+vWHbO2BX9am8i7ZxOt51EpphKoUtHL+wiehsIPSg8qlRXixd
5ALbAcUSl5l7Mt4hnjCWfxAadqknCLsV3GqgcJ6+uqexS3FN1x62o4Wje18/AAVvkU+SPdTnW6Xx
V+5iq0d07HFLhHc4FSV3LFH4Igb/NguW8sPYHqsOIMUQy1mOrrJBCA4KvcNGUFWZv/EUJpwouBRr
jxY/01uL06+rrMdXEqr0D59YC3ew1xIOUp9Vw8TX6iVQfCYf8k+NBYELhRqKNCqGppAJRZQlPuXw
uCfuK14X5rvCEWsH+uLkdo++K4IVIfShO7YLBXlstN37szd0oUWKRMmHqRV+4EuDiICtoZRDw6hf
tJImBQ/aWwkmN5mgqz/jLc1b2BrRN49+lCzmCAqYVBDgT54qEYIIfltya88n32Vwur3qyIHZhI9b
g15GmOsJkUXcdhjvrs4XJhrc9FqKi4eOWsXD3Eo6LJu1ys66i+9/S6+zgcaO4M91dg7MRr2Qfq4I
aXz4Pozt2o74vQdDSczGoV9OVHp4MhjKvFIQMVHx8Vo+DvEZodpX728W14EVk9RAqdkBzItdSsIa
yINOl0t2GQkegs5oRjOIpt5UZoI8hB+zgG4Lz68i/G4sadzg/gqDkSYyyXc3CnzBahBVncRixHtd
YsqsZkPxcTRmzaCopQaqz+2Oscv+aPJtJszYHBTRxXDsxDkQWLPH9eKZpmFFOB4sVUqfWyUnE21Y
I3g9DAUPeaVcIK1ssCQLSZutIVmHr5AVjq+bY7ZFgzg9uQ05OkM2LFQdGvvUT7XiQxmM1I9jvtdl
g8Gp3ywT1Oyx+ON/VvFZfRYoV4FFwcL82h9fyAFtHiEiSy9S9cHy9AxenelGTvO+U0QxKw4R1NB6
n/1i7/B4jvNEJLVRlY0sWQezsPVPEEH2TyViECT71OEjdlQ/W/1MyFLIYTmupPalD7YBgjeeAoP4
/Q9H8/oVUzS7HJh5BpoXZe0RCiJdhPVHWIUaC4rwIE1D0SOXrmBA2aZYWxMx6buKqRo8fSKuuv9O
/B3c+WC9gIAHeUVJ3bl3o3fVufa+10UhTtBqMRPizs2LtcQBSBTrUy7sm1K/FkiLFofmfOz0fm1W
9v/mPKhNzZJAbx2LPcDMV9KeR642X8EBdOf/hRcdoWpvAyCZdDlOQ++Ri/s3JyaAzoPt64keEM2/
GBWKUIjuy7uxUGNj2naqnBeuzhjcbF/OUwNY/CP5/ovbR/c1TXvbJPxDFo6EMj3DldKfY35dAxx8
K5fcQyXngwb3Umgct0+5uhVcviaevLGkAYWdA8Y5StPj9+DSB8E6WPYpnmneiaCZ+rBjVpXJrIH4
dLsNhf+5YQ4wL7jF7uYBOWMRS9yK7esJqEq2DUlfgR0TOMjXUcZ5+3jKBOI8L+G2aYWtTmep3a4h
9bc/H9NtPyy68Qx8/XWz6rsyaQED73w+ECyIhI5HvaLpxfYkS7DMM/6h7yzHqknJ05/uo+kGLUtY
w6pAX8Lx9+p6PsIHG2kwK1XxEM25EUTiNp8Y6wOo3VxTxUHpsdO6r/ZBUwT69zSfbUCRsIyAvLME
caNBATtePLu4k1ekgFTSZZq32g2qW7bZBU7ByFMU+5ovgskt4/YoldHH+h8I0ky3a5puFfOtB3mH
hhKgIs5jdy1nDEdsYjqBgVrflQDvfxBNn/I8A5MK+X1DQ3kdXYeqAo80xPCwZEgxbRDRpGpGqC6H
eY/yhggkjh43qZddWLYxtp/hPDSi9+8OKiN7nMJ+Hq2OyDkiVi5ibZnsyt4mDm+wSIyufKYLuzo8
nlfcxeN9XoMKKUvZdzTUmsKto4IACt/GZL6CkNh2oVLJiYZxdeJv3X9/zMB7TPH5zYC7hBQz6sKn
GVixm9JHLmwNxDe1HUCfaUl3SsqTeqNe5v6G2oFKPTLrKQMnafzfPcpPRAwPeDqATryQ7QP+Irmb
XoLfqFTn3CQY87vwSSpVfsbHZbvlG5IbWHRoQ/RPMJtgT21WadqLXxvlmkXrloJER+u5E3qDieTC
ceplHp3JNzUhcBNdnNZxCnJnl09xm28P9HNFGwwBH5vNtA73CVffK8fi0XSBLx5D3dPW4p9CHjJe
wUiLbjVSLd20ahd4LAEmJpiZP2+hdhdLQv58dQE1i2YtudKRDqoqTRX2LCDPVyizC/ulSMttFBc/
gxs0XDtcCX4J2Rs387gg8v3BCM5Fnj26of487kdry3Jz1DkwEuTH1Bsr5aK2GXpvHKQ3algGq+ha
9W3+r/XnAD6VNR/HhXbrOhyzas0sTnp6QJeXOCsdI2Pgvgqjqu9W2PqINphOLodo7exL2OEv8qTE
lfwQRv4vSGTfypOqVs10poILveumFEQfXFZzNeV4vxjC5W9YmI5PLG8sYWgKWVqYgRzRLAMsAkTG
oAJO+6E7a4Qbr+yQCY0Nw4jY2MZtpIEIMFI7JYlnQ0ELu2LhzJsxR28aSmUUR0mZcnOKiATARvUE
gdzgqF/2BN5okIKikrSvKFQ6N4qQAUo2DtiUrAF7aPUyfRq8lQi9XkVQ55aeM4bLvw39xRiRgmDV
p9yclugovnDj92cug/4zvqdc2rwg4DSzdsjIrJSLWT/8/2fskPvJK+17kOKhAXm/wTtm+HB4QSOw
IOYUpcoLuK41lQ33/ZcdcpFKKkArZNGy7zhLahpKbEcZYYJT1WUbrJ/JGfhjWghqBYYrKcH1YuZq
/XkGP1T7X1eaW6jfsMf5ylgEnSPYfBS/koOvyZzGMjKKz1+OKeV449trq/t0xY/yaxyfm8U+8SIt
edLX8Cw9AFdJcOc8zUZXx5PRy7GKcW1aJsFN8YDuTja+uOlmzh+VjGE/qNoBXgsLaSP3krEHzGwZ
yqNkM4EEPAFwq/D1Ul1dzGX2U2BSainkbQshtQMvaN2wAYlUaPF4W/N7T1+byz0insZrQTaCaZmU
618ijZhR4P+bCATgSDzPGmSw4Flff9aHbbEQteV4AvvFy728DBmpuqzRbMH5dGl+gaLqS4m7n/Ay
2MqCt1lsyK2xlyREP+qBs+4EuzMqrRTLAfLCSRWcjoQ/xqk44MF4TjHHyg7J8JdVtS5MkLe/+Pnt
qvIZ31idc/fS/Wk678NGKJbsgI9hXIrRcnYezCmdJf6SLsKC5kWUNGH0wDHQ4LVqgHF1bFVF1IVi
HNmIE4nG0xUlqrhsOiF2fdCz2iaKIXMNT1g4s8jst4RkAHkZmuP7qlc1KZ4YC/e8MKqIFuQUJxIg
S66K1YMPm7/cCw1hiBGRI35wVH/ioVKe5G7zGYlmTCmfn+PE8IcjLxtdhpF9SPMVJ+Pq0+Nv9qIo
e5R8JHpi2owdAZqDZ9SVpsqW90wuoOcZjSZIfvsl7RomyHzP+OfvUMXPm0+6KW1fKSQAOoDXfExy
/hPYdFNuWvJxM4tSFjX6xuU+rCYgxzo1a1arH+YZpexkx3bUGKFz9jRrss4C1YKWPkL0tgQ7pjaS
X5FX9spPfy4KMLsFWO0HWTE23sTT4buVq0xqDIl8emm4KRocrPR3fEF7OZCalWt70p9e33+PrjVG
D6BT40TRr7QG++oWsalyXGroO7OuETNCWyzFrxr4mHjFto3bG161OD6FGCU6X0LVHe8c1zeAiiOU
XOj3gF4wKYiXYRFGasnAhTWDTL30ExQ3bhIsIHW58zHW+dIwDfsa0XpWIfhk6CZ7LrSDZeUuXkz2
E7okvKZSTpwIMP1g/GkfkWsbH0a38vkhxLXnPyORwmSyD58W0Zgb+CeJATmQiSEPMb2wy1HGzjfj
WSaIR6Civ6fsPZq4hFVyp+hrjb0KDrccf1a8ef+lNH+R54xP+GaHpa5K5VLK37n5mx30Z+i8AuDU
rUoCm80YXcWLrwJEyidrLkvjdYcsW8XtdU8wOtmcgFQueQuNjrDA9RU6GlVC6BMghkak450Mo5ap
YTOSGtw//BII98KAw6yRGriOs+xCUSjuM4jmI2UA38WPL3yGs+hmxCYvoU9a45JJuZ3oHUCKxbWH
TegJbd1//cSuB57PRgTvWrdcGkGvYY1ZFcGOLzvWbyxL+sWOSkItw3hw+p38nsWcfQGuzCbMOT1z
O/VG0Em2zXExmcfQwSia0f7GdH/beTSGxZd96kuUcpUaSwqy8RMSL2Sj/8qMXhsTubiryT107HhB
0FC+ABrHdcJvZYI322pRMuyQJm6dkdMr7msvc1nT/xpb21QI/pXDFlxB/vM7pR5DR+bLuOuPG2ao
tLx4dHmZnt2CH0d1Lk9F9oM96qxLJOgxp+MwAv1OeBbFQdUIHDPI1Szk1w2VhZ2yxj8RHeyBE/DE
GpIBQPPllY3EC+LGLsFG7Y/fHrVEfIi4dPW+wCnBi9FqR+C39/A5ahvJWVAe4pkvWDSOoK9/dIu9
wgOPSQWSOAruHORbmrqOY4RMebS+D8bMK54mC+gzh3gqNA+YQK9vV3mN5d2JT2kyPt/4C2t2GJlm
2iEQ5VNQvj/V9XknigZTIEIV2AowCXW1AmCpYzPu7YYlKfYxsrQFxwqj65pr3dPfgSf+CgFaLr1A
jQz+FAradSt0iIxdrxrg3f4fmT4AkL5jYyq0YZ5n9mlxW8H5OkA06mmDWtDfe0453oxQC4syO635
PRpwL9XaYqGAZYz7HthDgHnGwchnRWOg904mJUCXwQKDwRwNfSUuSRf9TDhCqmtpvY8jp8oF2Dzx
LCXSgK/JVyfgyUBgHlyQnNvcvuuD8Ac/EVp2kfIwN4wyRgYLTUp7bTN/MG2sD8JboX353Z4b96lG
J0WHGTrHTzYyezVrb5UsmX01yTVzSn8bwgwWfU73tjyTSoGjDexg4kJe93q3ZbjwegehMgyOq0GY
BbwjbZvq9djnu5a5pnizwC/yIZbqLk01RC4zC+0Fd9IOxetzlZ8ad3akPCgtTouLD06Mu+RAs4EA
iS+xJv33oxNxaUtuuFTPVKU1Bt9QZOW88AbH0I2CuBw0deCw5dUtb6XTKjvrXKWV6Vn7mXANhsE9
96cexskWgHTFB194rPX0Hh/oNiDGseZCxLl9NxRataTZJBDLwik09hmmrc3wyxNmBZJHSvtRn/H1
zXz5Fgvla9iXWejwDX3+vDSxds4frwOZ/yyShxaWTNJVT2EKzShZKM9T7vXELHwdZ+9KH9AnfViz
O2/zImYdF4yrWL6mb8MCX/uYOU8291LvUazutfhj4HHPaN/K20V1cWHdg9cpbZ/6NiZWWgEVzPF/
jBchNJ5mDgbm5Mr0u4JORRnqbC5OdrMsu3ZrVLJmQ7d/wrDgdo+lYz28y9ymbs+OpCKEZ1XDH8/u
zl3BDt9NdW0hBvQrzy4lSDvKawuY/g3AM7miYi8SUKkCLCbPNL+MT1TTiTcBQKHt58Od0jkdrOUI
7U8opBO8n61E79q5hYBcR6UNkyqlRjG+8BZUkVZSUe9YG1keBtsCstzIben9oybn7MVvnIJW8YoB
zZg9DVIAs2rNxMLMxCg+qmtycoi4z2b5g0eyqtRGCr8Yq8A2y9sI3sQy9UoWDqEGjWa3w4hZouWT
aOFLKWGycJtd40TTfkc3vACstf9hxFfMWslRK3UoPmXuIA82kKvsupsJezOVaoxi7rALKaadYNUO
bVKSV8SZVVSuGaUa8gJzk9KAizgCfOtPpiqp3rgsTpb1az/F1sACeXwGFyazPy78pLsfmEVZDgfh
+A2gJQ3Aw1kqk6p+6Pjc71KrnHebbDzTVUvZRO420lKotnEdNaqVssIVDVSe22ZQDgEUeW3CH2P1
4Xu9qAg74D3OpW/+eIMv8U7fHltmgcIiZzHgnOlkcfVUflNhOmliIq8Gn4BAzA4Lz8dctdmFzFZz
8yYkTnJ4Ow1tUWs5hIvDqkhWXNggXYbbYCcPK63BfyNSaYvSpsTP70G0yeOgC+m+2YwA9zu/WDsk
VJgxTPNBDJswoQNWSbkjBfYZfaCOwsuhjH3FARn6lwwnMwPx8rC02uaLKlDj2S29dQslYLNsr9ij
5T3miX37cF+vuRqda88/96mCO149TM17WEoXpZ5dXOWvZ8DpFmfPk22XLNnlBesuGKv4NX+0SU+r
8J8N6tlzMCTQ9Rik9a8nxRA0AA1+p1Uaux5nPVz9xse0BMLxxD5ki9XSEwF6YJXSzFUGgN1eUnFq
cBVy1R8DwgKhXP5KvkUeFCMxAQq6ehkbqoMKi1Y2J5k0/BL9xfkt1+5qPBiwX5rRHVX16YAEZjsA
MO4CZsgE2ib1Jaoux9+DI3exhbzr3iCxXIqO1DTEwZcw+SmnF2BQUMephpmBN+j/xbRjpByLd7lf
gfySFS99le98BcitzZsnv+hylWjPk6Ey5+3UB/hgkFyJ05W7Jhjhh4+HQtjKQeX1eKPVaSsbxFRp
Amkf8V046oN+btcfKlsX+QgOE0MjcjDz72GBViqruXGvwxiTXZG6JtgwPh6vRYyV70hn84Ool9r1
YcN2lAXvkDEVbl3yqryvElUPSzDPn5BkTDJnB4mc+fBW3drutytcYc6a/Doa6wKw9ZaeH/NvtrAT
zvKrf+k21p5j2EeoZQTIN3SG4x9nOVF7OSJP0vM9UWUsudCCL74asspGlMUNlGr5DVUvjHV/ity3
btt0ma9UsS3iF4x9Hm8+5GlFi3rFD8TVZGaXTp6FzOjtVd+abmSmimFWBB0dJVwtVqylhDQgHXSj
0uL0wlhYfXsynGBRTxEW9uuaiA9Fsj8rqIwO4WMwVGSrh3LRmMmVKU8hRhCCyHnvYZ+fN4H/lULx
9G/mcTTIaFHhglBtjTjBbMghpQ1BuUVpP3+JBFOBGKiaM7HR32uvbZ1G8LZDfsI30BhtqDWStK43
VrFW96ncrOVo/QDgRBN9VxjNr4kn0Q+lrA6q8ABQCFd6sXiej15a/upLNeN8W++0/eLhsSoL4QNV
J0Af0K0UBbtb4ScffPwf46eRs5TgXWtr+0HIWSqdO6fU18sAD7cJSXtgANDyGHAW9ZLaH9F7eaP7
XAaSpRyVYeaTbvVtFKidrcE+zz08XE2iJvGydKuomGc0xCUitEynf95zAqOUJJ1RP+5uXxlpZQR0
ObYH+FwbWUu4yhol1YzKcgSDjFqxf9jYdTP3aMqVUVhBwVkMtwrPQ9cntQKFmZf+u9Q/MMbjEamz
5yJdIFhpP/EDI4iyhp/MGBhtmSi7CkAcQxYYys/L7/bwqD8YeULcH0ZGYLkiQMpreWAk7sPsXZJ9
uh8S7lyRkp8SIbCQ4VsrRqk0q7+Zt2VvgvfPkB64yLUz6ZeUGd1t+ps9y8c2Ic5wQtpmkBDbsqpt
3IZ1cDJNqCd/yfKDV8NbKY6zr89xl1eHcJPJfWeiB0sFiw1X0waNHPWsfFzcxwEncSEzbh7AOdzA
WQevne0XtxbQu/KGCYHYl5KnXXnr1lUbL8yJqBPAfL88PFY2kBfNmWuzRRyu9uUR0xA2GcrB6lUg
pye+N/ORzHM/IXd1S7qKl3YOiLpmSwGX4iMkTVx0kqXKcwwY47Qen/2ez2X2UJ8rRkxWya//6owZ
c4YGIoRfjjCXAMi9GmANetn6UHRaehm8HL+knNfbOhC0pyB9R7417ld82xAfJvfcVf8bgPd9lV0j
djajoySbZUoCsv74D4hlBX/NR2k+RKmU9KRR7qIld4pm4xc+TXL0YZi/l9q7T65ge9WbE93X4KTD
CZD8UbiGHd/DG1PaavpoBBfixVago2DuIc3r2JMwGzHNC98ArTdtWqeIrHwnIBEAZTsjPNyFosyH
uZ4yrF0omS2+6ygMDk3oUVbDLtTlSw+2sSa71tNyNsW9Uzilj+lph6KosIq6ocWEkzUb6d3AnSPY
L1wtvLHm2duoaBJMacHAcEwh+l54xPRgk6aJ6/Gju1IJtCZULxsllKpC0xPluEP8iYd1lsd+Rhn3
3fQsVulMc5Po5Ir8DtPs643r33sQq8JsKMFUUC7o4HLiyOWymdtjMZ6i2XgePVAM9skxWj9UCOuI
CHAVl9gr3T9i+EqllV0gAoLU71gXEw8RUoWWMNkQETgCLJR2ZI8TOXJxrngON+yXAnlrkdsTdEK4
rPkQ15/7uqLH1hrIen2hIJNFoivMuWumxX5P7RppnsUuaE3Jx0YGV1WBkiZR6DXz29zwSuqfFfUB
zHcJPAiHItmhQDHmzltB0bpe1f70z8zAjcNoqwBFfOMHowax0FL/Ckq1G7wPxucbyGTNNqF7A3nk
5nkrMSgdOZ0bKehoRodqiW9vKmDJOc4kvgoMvXbXBridPbfSZWng+vvAsp8+I9u22/7bAW5RW6Yq
1B8xo/g2Qoxga0KBtmCJfhBD7Q+67sgsU+FT+aYRxzHSCDl+eEgdK/CBWV5QlLYeZ1N1Z6PWDIa8
0puoHFXHdYdTRzC2ghT14EjWNnOtQjJ6+zacScbcV1RdlIi/FOBvrp6x12ATxuAvRH/01GQndrcp
a2vWVu0+8R61GcQzsptW8qINznqTYiS19/GeZvugIyeMTv43wLT0orKeLUs9eDYR7XeRmC2tfMbk
DobgbjsA1chPvUvr2CioaUJmTS3rhJ+UftKNVo5J4y5ixYxI7Mm8ee5ErpI+gcJJf1tR2CP1S9dC
512kOQYD+rFozx0527zn0r6W0PYC8ZVSbnY+3LOSsNGS3ooInGk1D9X5lxV0f6Dckmgyp6uTATSq
pKE3J3pVWM6j4ZumlHidk/KGkw1tXUiCe5hqLMdd2zff0jaS7Z8QcRUc5sbxNH1TPhNTZj0O7X5g
sHy1jrI+EhecWp3Hj1w8n0m3d1XpKLZ4TbKEs8yi6WXywEO8PCVOorSOPB3dQa9be5q4Y38xkELJ
z8HO8IVAhT08zNd0jGhfytRnQcVfX8VIc+5fNGawzj2xwFS2qlNE8RamzOprjC1tzkpzotu+lPjo
B2Lz7p2nshRcIvtVNorFl4Ccwa74ClTVxzLfplMyrkzWbL+tj0BXwVW5kwrGizn0AQl9IGnNsVhc
B6jLd3dgs5u4UqVnNswSGc2YY7YLEHHkYKtNZuFtvtKrLJSesaI3haoelrWJxaQ9sFEoOuK8DHHj
WCw2Q/Ezob1/OtltQIy2cbztBr3Gv9nDCr5v+7w4F3cgu81upafJ/Yf8X9A2Bs3jmuFtUOpRK3+N
nt0xzlkh4R/xm29137JRdODiZCRONHk70cb8fJyRUNvLEst3ynjiopCvm7mW97UZ/MJgGLEH9vw0
9k4bJJoikGIpo5jm611nk72wt/NvaMnoOgKeN1FwkBr9gzU0fBJBIYi9hlizrWIvZlQo7CIw6WpN
OBiDLHNksD51LXAeYKC2WTHBK1Pq1AoUDzFjONI7ezpKmVPDC01pFwei2svLeDcTfoL7tth0pjH0
sB+pCDyU+s5kB3Z3eKn9got9nKB0Fyr+J8MAbg8JJGsGSE0YUNTxLmTqI2l252ADZDXClrx1anLB
MP4EYEGcCEgcuizF7ucwjUdvMwzUkHymBQW48FAp2gYb33YEPyTWFls60sAcYJnDkH3vSwlgUS1k
jh62PbZ3L9kBsUiP1TYe4uY7+bT3pd4CjwoLICFnVsnj08TWx+sV26PUPScjOO5o7sBY96bomgUC
ruJ6g7RgTD9x9zuf68GYTz/wTX1EYKnjJLL+GbeSKt/3bW2jJEt9dvtNLv+dzA19fzKjjuEHFoOe
GzMDNlgFEiBWMnwvVqNMjcpmY8brZpS8W5W6Moon9FPrsQDRJIcX6YSrb5LWULaNd7sl/TY2c65/
1RMg+NjIXAB0RqTHD8NJodWqJ1NDsHsHly6cv3lyJPw93rnQ2sSusc5kD4LvLqWzGNdWIWacLkyy
yRNiy0zc1nIdIRIsBPNnm3CHdVdpxCuvjJKBtaLEqaJW2o2I8rnR9jxw1r5cc80Euo/DNMRlFIlt
RNf36lMIbXAvlDSQesl8ZQlb3yjI/sdzTMVLSZpGeE79bJ4nIL+I8WW/kwglqRXgtTPdpIoxzxhx
w4m/VmaEsKO5KAC6tkJS2gWi1aNJBtUzJTICKTXrEhmSvvn107HKzEUzAVV/hrhpEbRjzASJb/Ka
4wCSROQzNnYoSbCPVhHKqL3pDb29oWCnnTlrqGUwksPq/BtAN8KY0G3DwWyBRP/3EtM1/gkAUTt3
IqqObRps1mtfbq/eZjxFkiUP11ZI3fgZkQeHigRvdX4AGBPExRML1wY7QfFN3Ym4BCedhqymyGOd
sjKwQ7xNxc6asrQmn8Fahi1j3wuGjxs+xMOoxGKvh2DyjrCypXdrT264gX7+Y5pGWodbM2AdA9ko
fXD7YfZ3X4ERH4FWDZzvfd+h+xbp/l3/YLlo4w0tlRQc81AbM+qfeBbGNcygakkj9nyrVZU8LrJo
CryVJGyugl2U/qVNjkglgevGgni2/WTQvrrSk2nXUO9GKKI73QJuHTweBcaxx2SkrHGkdWgV+LFv
uubv/cKGnWG1ijIejdVEssPavUfMDeKPRoP7w2cuUdCLQpHpQIYjL9UHeGR6sq40w1P0VK8enBzX
b4EJcxzEzbVrXMDPG4yFG3yjdBg5feiLeZlmEHI07pJ6B0SjOMt1C2Zy3Yq7eN4oSu4+IU8KxZ1K
FAr/ogyyZpl/i2bQTE6pjnL7Hg733BkbisMOyEceTBLd+ikwz39VSH/l4TyfvFHZO6SjO+v4fHQU
l9wKJfz9j8H+Xjutg3hHdMrhROwOZmvRMo2bteNTwpVyi6wZ/t9l1hgMkrRAqod7p6Bym3pZecBM
JtOIqcZCD5QGZWMR4pLkKzRrK3s6T2OOYlLocKyqC2D7mn+gL96/bZyKvpLyymtsFt7UAJLNiWAB
3eVWym0jGtqYALdrVIhvOCqR4WVNaecXSuJsliI50Ptq9drqwU5D8d4QsrDsEKNcVlYIbCVYwvfG
jgpBBaRC4K2WT0tHuYwhmPo6BzoxJpVt7yUU/nBEPsxKRmOtGb4KXKknjt07KLxnlIbY+Rd61E1u
aRCSU4Fv/UWoSbC/Iq6w+4cqEc7WQ6SO7duD8K4EMBnZF/9gBXdBF2ZysF4do8dE0eDOILez3fGO
NS9bSkUOhrU+njLhZf9gmHL+ptwTzYY2AD9s6rsN/nGsZ0jgeRcQdk4cyhn3iwF7EXqewkWuvFP1
kzKyqxJBQDD86CbF1EUcEhZCvbIYz1cEeX4qQEvFZl/QRMjqLorzkrjt3e7bqj4p+fSJwnfAmTg3
7rHT1UIJO4FSCDq8s7ZsyR7u0wTQHoSe3JC4qimI8ySqeutgYK1R5Fdc/QVjq3V5JTodhqFyx43b
+Pwv2tE7pReTj8EmgV4abmlQ6O++Zvh0qettkvHK9GWengdOuVW942jM9lfxhASDiI3h0kBaYdA3
alQm7lo4AcQU5ctjn4LqcDiCyaA3R8rHkgpRsGJ6OYW0YKp/6IcFpNKfB/5jbHshSJFH6qhgwsnc
/OuqriQ7zmdbudlIta5+UrtUs5OXsUdxqfGc4+I4SW2gd50sunczUDvttDhVg8bheYD+BynwaOp8
eUNExsLoA+Mf9TxK+g8tVyntzeQWVTnm/RhPIntqSwhDE1u+Ak06kvuY1UZ1pDPutbVyOxaHqBQ6
LtzELZQxwgrRzeS40TdMaD2JWi41J6bsCJ0ElUo4q/N0T6wUN+1CrTUPGHLSIDAt5/0Z+01B5kUR
nByjwBHtS9SKupsdBWlVyca4wXObJMTO+zgtMEWVfF/zeuDP6ALZ0rDpX1tT2uDazN9XuCmRORzy
vp5oPeKV/MFCYWPgnLXDxCzt7oWHy3nhTXtVWJdcm3IHrfq7XoVNkIqQfr1UgfcgmsY74wqWiZ8g
I7A+ukV8rRYwcrBRY/k+N8PU2VnCFTXcFcdo5KR5xf7NfLGVFdbsAzzmtBj3ua9hvGh9vbx0Z3eg
AljG1clUH+SL7yyMMxUkjGqK6R+1A4ga5PWohm9KWKAgX3uv+A6/l+EdeWRkHbdUfrbl/dqmKKto
70wu51jyI75k8AmYur62R59vp96F3d9zuLpMzw2Az7klIEVIXWigJzaD1rbAAN6m3BWcLGrcznk6
2/4TyGorznc+eW4MPTNITrr5O/cOdLH9tAKnwQ3n8dTGvXDcAwFpO6kcOgMdNizhwXkMPy3HnvKb
GKiuc0vZ7boim/nEZ097D4kfPqU6Og7qAgPG6VGJdI7Xdf2JYNdvGadHnsO3mNWg5sP59vg6uV3d
hdUA0KYqJGyHLfGpeHuIseAQUlwskkGl/HjZGo9M6GnA0W0nWKBxLbc8OpUAhiigeJbhTY48z3Hi
jN5jVg20rj2kWMdOBUgPi9NXg80BodNVGigwQ1vwY/pKVkzCodB3zSI+hPcgq2i1h+zFv+f4ZX/T
e8KaEh7MUecBBR8UF1ArhIQe8XZsOD0ZM4JdQrLqr8acpDTPLzRF+FkSkItVjVbWLeO7oXBY/zDR
BgMCl4Qw4bRyG0pe9GfDmHdtlr5/D8OMvKzduHMHsHGnpEA4Zpt87jWaEJ4JZylWg1miYxAAv4pY
S6mj1WNKOJ1eAJAgcArtzTz4rJe6fhnY/wH9HA2MLM7fBeVVFSEjK8Z0Z/apIdiQXvJq31s3qFoP
hSOCHHawFeJg+GH/xfVlZkv4ILLKmC3U+a3BOUvTVUkKowbCGLiPNtrUi7fnwxclnFdH1Rt8Cm/T
fv0zGJVvbgigJTgaHyd7rBdepXmsaIU6mAQzP7xsehlkv3VBhZ2MhrFEteZqMUFNsxnL2p9r231x
s0ReiPG6oX8Rc7tQHJ3lviGMLiknyVKSX6IAUEtQTTrWcybEjxklBX7se6wuzo1h+oYDYINurDuN
XXy6HwFVbVol5o6wvzXaMz9e3J+gxR2pRsPqxnSJgRfU8fApCxAjdL1txms91fuFc3vbZFW/kQdw
HjwWV4kwOO7bbrr/NukwCBt1VaS/tG6fRdpqEpbYoTE7EI536IwNSuQtY2D/E5f7SvZ17UN3V4QR
dZny5hkaWHpN8/We4eib/0aWJKy4EnwKwNMthhCiJ8ftmcI3uQ7hiiT9T5/36FwAx7neiYEh7kcH
LO0gmEk3BGl2CnkzWYcsEWDwEn0J/gE9hLH+V935iE9MudkeKNtyqBFzwTBVTDwhD5aMPpgMdqo8
bhRiWA3yMUT/DP726ewylYCnTEknF3BnbPSmblmqdQDMpAAKJAp8ezhGiXoNJUVA5E89+x2jX7GB
ok0+q85/hluTrUouDhwvrKa+jLysPWdjWohtOEBfuPF6PHN1L9NOe+17f9XMkX7dMs5WcKTsmiBE
MueTXoIOje7heI7nqNrbtgGuCC8XHRgowZ0QTJZ6dzG9UmwkowsBGICYSRz0z56uCin013Tm/P4J
MTmFKC9WngYWNul1XdwhEKUz1Td94p4OARkk7fUXAJ7Mjrt9bf8k+jC+0P2MiefRZVFJIB2QhyBl
ivNw9+e2u3ACbhe/Z6YzorlzsNP+faU4H7f4PurU9a9nj7031G/e+zrcckvwmhya7FXIdYMTEC+q
E5ZB3ZHzMLWT6C0m/h12vGJoEoq8HYh8/9n9ZqVX6OF641JTnI2OnEjqVOb2JtZuCfSNA9vRWm1x
Yiv50iVzi/NtZ8a0D1VKnVtkKaYQ4izd2bil7EH7NIFYSsFCueLY7ufsba2XUFLinlv4K3jR1l86
GArcPIt7TYxqg01hjv+2pWzOULzjbrbL4KLLy3s74s0qvhERr2yzgX9OhXNtmUJg89uoE7qWdfDr
WtkkLb8DuSbyEuLS8KVREU+bYgfrtFI79jqrftwSjz2+MIzyKsn4yv8oPI7Mxyvw2gVFAOrd8DrU
R+VVIurhNg6+nJwxIuUU5Nh5pSc7lKbp455Zq4n70hQKKPEm5fFvepMxpFYS6RtHOVVWwSdncrJ2
X14dwpU/BEVqPStqzuhRuVlYPHJREAwRAswp06T+nX3XBg67alo8BczTip62k5fFeUi3O5GB2dtC
lHmpEvKturfhRcVVqymRyxleZfwrL73ZyCADS3CZue9ZxZ7l4+ActBcQ5hrKsW3B+rKrbD7zNniv
hC/0k8gPd4PRFeCSfSyM1IXB6soh4wxhAQ6IsJ22li31/CLZk5tm/9U0jKYz5AxpSm7lJg8lMYy2
aFNVrzDVKCtPpPFnufni624coLykKF2LVdkako2cwnlnbcbbNpc2pm7n/O8UQXxczq1Mh1NwiZwH
p3lsFxxL0PVFd7dd+mCyWYIE/aqXciwugm2QdrpoEgCoTtw8zuR7vRW6HZld9fbEdu6zPIlLvgLN
BjWq2fteGGL9mSN5u3B8DtXSH3gpnXJ1ULZklfZUVGid9qrtzRqBf3Q0pEElrftIBAQG+ksHHJ61
b6x32RH02SY/JfzK+zMBjMw3rOCgqio2HD3sRsz9q7pMYpmCSgLQSu06vuuSoixGZ3mlHDmuhbvS
1BkW1SHuFjo0a3Yovec6G7c+hqinpmTMdHiHddSY2V+qq6gMK241bSa7/2b8zJzIQ/HNoUWjV72p
HvLt5yM8CRASVVuF5aJPzCTtppYqjjt+xQdn0Ec7G6DjAtuMNYYq8s5Y+gUORwWOotFstutlsQk2
kq94hxLmgF6GFv8Hrmgdr2BSgd3ObALR4fS0b5+8sEFie4VJCanKc3wVjuIffjkZSeSUBTh+zbPT
eJ6WupFknbRhbXlA2W7q+v3pXMmqpZsFU7/xty4Ndx3bBhoqaAz9eHsodr9jApUAGD9VGxUsz7kB
s4Ikd9IdIqRkI6KLfOikGSYuCnkH4n5ttK5mKyDww2fZruqeg3wY7c4o91wPE7dicoxUz5u2CeSA
U449eBxxBauGVFwzaEVCCDLVdyNuCK8BxG47tfLeY+cnq97EWbaeUKxi9GlrOM2O3SVzmUjpMzLU
kTv7wAc13le2+IAveq788mnNHU0ExqjClPF2RXNXEC2E9JeOkrZ1VAHxyo2vdatee31XRJUXE2ta
8Bwy+2TXqdVQS4KOnxk1GoKjueGOjffTtCgYykCsNV7ejlLAHh/h5zBWl0fRRBO1CbPNrtlCe+Fw
bh12Gnc/d3nsrP/yUKzI/hIlNVwy0QJZ2EtB7cMBZRqfcRjWDuz8YAfrL8fPosQZ/6h83TroIhPp
uGoRF4UkaOjZr8rDCiOpahHSu9l7/onastKT+B7RAXB+ejPB7fzeNajWItEcyUzmgsg/bTL4Izm3
A9g7V0w3AjXqgq6sE43DZDljD8CWw7THv4Q52YKL1erxQGCJl8mJauDxXHE1mIG47qor1kMzYLtW
IqK7QyuntP0yIoiyBY4Ql7kfb1s+r8nSX77p5I/Xakg5axbAMFnOu+rNPDPmbWK3EPVj4jX4qtbN
jYwSigf+I4QnHHMg6pAQqQPA4y/yKPEKgHmey3LFnRTGsvwsfrUrpqiNOJjKv5tIV02ZIr0XKerC
Xv8zyEnywoafZCOppXZGy7Kr+z98QG/c9V/DmN2vKtqZYPhxP46Q9y1aP+wvjc5gO+OLRoWjvALi
S+IuM9GNIfQ9tggzuZ+8iMWbEUmZj4junqThP11bHLBaTGujA6Ar+dtQxw2tgEHu9L3d/0p8DvV3
2y5DU+ExLU5BvAYreMfbJZNEGTmzugqnVg2RMqdNpFiZ6Ol3bqYfmdGJWUTtjlHY//5+iNFiLb1B
fItet5bcBx7Ohx+jbnDQChLLvTPYC0emdbj/KLk6YycAMASmTp5v2hJaAWFwr//vkS+Pv45O4Qu4
TAZNukuRJ63gebBrxmTkBJQ+8mKKZqu4LdGuZpV+jzJHrNZA9766FDnYVyjG2HwHoMdVdT5TXPOw
5JBZDkQ+kIEjtKu9lRGHNcRLmcbK5N9EUxE5EfJgSr0Y++vw9BgW7MCeRRZ8Wa+LsUfrGk3vBjFd
lHVw54ysI4/ejm3IX+EBRhBp2P9+TBd2qK4YNh1USVrLpFN8qegPwReC44muVGO72XdQ+MHKKfwK
8oxOS/3i+GfakucjQJC78/L4++PYH/RPphDfuOvKlAq8z87GWT23543gpWVqSYUYnfVZGM4eMJwy
DnyUfj5Jl9U6/iZaY6AG+JFX27P2YpRkXORv0gR6ZIGek4zNlAN1x0ekgZyYHk5XrOXMOfktI4A4
rfeVwoE+r8Yi/UsMYOOdk6xBloSTVZkrqqWS28ANSBnxXEeHyY/T0atkXr9deQBaHUZJ6/mExHgI
YRco2MWlqfT9kobo80VCm7efYEVDrd09Y5b/Rm+4QfH7Lw3APVtDKVu42D+QJg4LLRIkvqVdWYuh
jIHgZKVZx1V6HJ6YrZdCpbzrtqaeBpHbMaOWl74GDBfEoym055UPiJW5ZAzu+uTxHik9a7R38S65
zxpqw34zszjZ4pwL7H2DHMNZBGN9bQhN12rY2ooqHJ1tyTXTsRrsUmlgFgAEkK6yLbdS+/QN81Sq
zorthpQ857A/mRY6HEopMQtUdSijn+Q0FKzkW6amO4VC13lj6GT59y7p1i507RybeMn26QRpvZZX
QAv13ly2fWpCjc0rimjEbm9cPPr1BX/gIvmmQKe5kPmk4H2AiE+blB48uUYD31FJeR9rJpkQtePA
hOHjT1paGhFIYD1clO40lorxXr6sFU7DBsqiquGlBH+YJZKMHuzZzsV974EsosuC/ze6hleD5oR/
O3z4lQutvXP/BA+XNjccZ5k62qsjGWgpXzL4ITe8cArYPbfQ2+atfF/dq+vf4UqKXD6Me/ZGv6D9
pJzQZb6HDjystrPrDgvoyVyeWNL1VJOdpQh5eB61ZTjejhIHOKBld+huZcjGdhBfykx5h5cEfez5
MxCF6prRd3ociuTOChMt2T1H9wiY1BjsC23UyNYu1nQFLis+Ci7IIC1moF1HyuZIbNXrGz5q+u0M
X3MHHK8z+I8sJkFvfGUVaaRxytttnWtpNOMJkuSaQE6/WG4I6Fd7REg0nvSjPJKrcCX4hE+UZgCT
fIm/O3LSJBNqlOk8PlrxtS2Uj1iHf9oGgGvvBlybG3rj0wmjqmVSk4c1nBBL1h29be2VwUHZ8he3
geFfezK5Ulp9FLDU/bDE6pgOaDXAr8yzbqX6cHRTO0HWY1POiFp/EyogbE4QvvCnhbvGryTHLFc4
DZpcs7hNGaMl4QfC5uILCWZs+L86bdL3QCADecOYPOhICXZnfcAJnB1AZ9bgWvcnDE6zuvLu/uNa
6gWd2a13EOEdb11Uo0g/asu2bqXg0vezT8YbSOlw+2qVMMV7gkXr68EIadxfoI7SFIfzlPtIiP70
hzGnSsN25G4/TGD17f2aVSoHztT4w6BalIHnH+eacoB7K5gv39P/t8k22qbg+363h0vS7xf+FuxD
Su0a9tAChM4PG7t1ae2fd8hN20X91RNizj5NIQbw+5SkfowuOR2Pxv0riabSKs3/dmAiI47O/ttH
pf9cbQtZLuH82mBRr8JPDidOTB9mqhgpqGUEL+zsCUKVmSqkEByeJAVOM1zB3cki7C56x/bVZ2as
uHL6Xm9bUesJWqqQI0/hbwpdR+7zUQTdntpIEEFFgWZMV44c1uU9EBBUXUS0XWPYHi1zpaj1C4Ah
fk6YcxfW2S3l2WRdAyWzOBVWMWnDSOF22P0DU2UzzvOr8FGLrLL3x/Jvg4hcAdMFuSZUoRqgPVs0
niCouR4aREgoS4ivF1l5Imq17JcjpfidjjHGnnsq9N/3tKLLtobjN7sRMBBbU719X7rGqA2CNc1w
xfA+nr8nwvdk+Cme5U90vh3zK88lywcYTynYtyFBmouD9EPdQNrim1J5yhmUrD6SWr6bQ3Ecrr92
7/PLyeh7l45iGUKpUccnWrP9nlN2jQwfBeCA2TMEXRLUqMtk0yjjd1usj8VLI+yuthIQEVhE9hri
DawBP67ydBd0Thjrdosh2Pgncnicz8QuPYgQTlHLKoBSATpCHwEIMXXLCU0ZkJtrjqnZRA9q0amQ
bZJLnnLU/CCNiarA7aRpV7H7/VBHdaIq4bWoskZOVjk3Rd9XgzyZculeGnzPFQ4+UMtGPQrXtbHQ
KgyQuqGTsm/x9adaL/Qmvla9/rDgQ6JuKcILPRKdzD+rmtr/EAgEtYD6XopdHwmssJbdxPW9VE0o
JQbtXIiYVHB3PRp/5+50nYah4CjCxuHqQQCKbEJ+PEOA8mzEdarLpMFi2R5lRPXEynOsvWnpU58q
g68d4bbojjeZyeaS1huzrf7n7j1VLx22ToLjOmmdT13oJxdmZ23bvT8Rlbh39Zr7p9OvmIT/wGAb
XUz4aJj9XPSxFJqfPr4XvXykeHz+Lf3wEZiFS88etW/138E9gQhJhRBF84ME6NjElINrKpDpf/7Z
drA0ycWigEUV4hTWDFJY0YvmZlsZLddUa/GqQYpmtt7CX+i8FD3d8r11kMF3TabYQKSEQ83Hi3Lm
lWsloG6JCd8vXR4emSZmRO/0BKKkM5I5jWuhpRkBNlLkHAt1sKtpF7nOnBQPRIAs7uCK2xBdTrlv
Ud8Z1n85nmLEd9v1q+zsHj8I9rHYRhUNDcBDyrWSO7xQPFYmLz2OSA0InvFzAiCBr00EKKY10gS9
pYFOpGy2R4Khovc+PdPZkv7c8J2963V+UTUhzYpGfh8kYHyRFF5Wstr2sI5zNMHNspU9/pi7Mz3F
gd3Qhm8qQjQWeY6GONMx2VHsakZFC2s9fFZmO754Oxk09M/y4vQPXFV7UJxJ6cwQPKyNPqkx9UJk
pXJV1ZTQ4wHgN4+GDGhu2cUkqYACUPr3o0ASyM2NDUQ7eaX4WSu8UKCY4UrdbNGx3LSjsE2gWFto
i7agXM4IUILOgPdzfzzgH4hlLC2UIagjpMhmL/hu1uhXsIYBQwDcHvsZAaOpT0+4eFWttD3Fgp/n
Z/eikM3EJ2dp+YuL6dxwXin9hvk4VL+0bnbNFoH7fdwLObfCo4T/FmfDseDPmWcQtnmSxCuAGtdW
8BNn7+hZF+SqSOwgIBfX9AI+2sEBIumLNTRB/lBI6M1j5qSY1pGyI4pC35PFvf7g5VQ09Zjv3upX
Y4UnVj2nS1M4WVU7QHNVS+YmfcV//oPMoZqxaG4B9BwVTsTyBp4/K0lPw6WlcRedAjGa2X78MMRv
S0lt23yN62VD7Txdumb23sHZCGQC5Yp+MKWQwel/78tRWuEHpW6JsgNSvTF1CK88ETqvB4atcn+b
dIQJGzcnVy2/93vGFEA5dVTiCi/0PTkXIvMXvGk9gOhwIMB70zlqJm8MLpdu8O5ofZxkNlZGzClU
oWeECUKLNHdc9qyymE8PH//ZRoohvk4hV24+1Mr15D3L4bgklsfqmTF0EdAoiSVcZYKDQSvE1lNy
ZWXpXgebVt24VVUU2Hq3PYzliTdYRgMmFh3wjCVKO2jI5QEXwIw8mNPn2OTHcd9N5szZZezCJoDu
FpuJJM1/5g4GN3DCImabRFHnLx4Kx4G5W01MaQbSQLhSyaGiCdSehkS9QV70Qpt7/pHftdq98X5x
PpgnA+r77lQYC/PlVHFQ9ICtOCH5TtLeuND58sZvWuw9bjfj4cY1qGUQnZbNGszdrkAuPUVs4nUL
BRuPCS0sKgm/OLxjjinP8MqzTRtduqfCzsBBosERwjQxYJziPfmt9uAJqsio2X4pe+/URqkW911N
0qHea76ATyPRtlyn+S3QW3XOZ5h/9XuWW7f+WtmA2RE/++OazVVBhQv9p0QqJrDEQB9kyXcHxjij
+xNo96JpNYGyyvdY03JSrwqqWS9wDZIzkEwqhmyO6ihRJhrgUh4bWqeFxzA8oa8ONMMrIYEfy7hc
YbKGgvpVFXow2SBuLSFLydemvcE4hupFxswOEkGDzmJEJaqZSXzzZNIRjxBpcxPDVHlPvl36OekY
+BDE99XeDv3yQkqwPhrE2y4z/rHNjJ7RIPFMt1lshQmJJYGD3QyvDtGBryJ1/Mug0c22iV6yMa9l
ZdH5Sy/n6WyZxQJjEHdyGAAm1tPu2bgL2eJ45HwJn9BASL5JxbWcH2mSZ3qPC/V5vktXTmedHppK
oO5t8caXtwxyvxZBrt21yY1J6QskZ7bvhlkB0p0mbAm1GKf2ovegyFyjA5BuvC/Tjap8rWiteSP1
8hrfHJEmspblstBC1PUOHHfcdg0toad8B/slrAjgqEZG6PximXM8B6C3aA4B4dZgsERyL6WURs8o
NgopvwDPkOU/EmArVXpdK8Muw4JFPO7HJr5yjkoQCHEypE2iU2s13TTxa4plxllTPvqxnhfuXlhp
ESpHCRpmy+k5VKPMIkXNH05TGHUKybMH/4mu0hp5rIWtBWv3qnYls71Jo+w44tjeL4Y6+nh4iABR
+MfrOXoDJFwb1X5sn0ZzpssDrnZY+o/cMM1OgmZ4kfERiVWXGVZwRE8UXTV63lEdQrl2lOvx8EKI
heZ1lW6WPXJTJmLt8X8hFW3rlvsFy7KBp/+5D9U+9oGjoZE3Y9RTCJk9ISTAXKdNgW0zvpPP9jrz
POmC/+TLP31PRB6vEb6nIk8IIJ0OVreO2oXj4plDCwWvwSPNQtbZ9pfQJE5uO/g/hnPqNcEMxQGS
xxUkawDmQQBa4YkwPWCfHHKhelgK2y3H1OWGDcFkAOgIzG8K3gDTLqZhsfRGe966NT5uWCvpb2EX
Qw+X51oyBosmlSn0BUg7U2RHwS1GkjCH+Twnkxn6xCf0ax6VKEGK8R61Wqw3cOndIl7YGuOXWkP5
p1ZgZtfJ3gadlzQUXIZGOAwaQq+EHYxGP41+YWcNXMHdVobHmvMhgXPGEIGLVyfqJWN+CbnKzSPa
MAUm1r6/vwLiAJuiA6YB8uc2JP3B2lbRr1rcmw1ClyiaXasWREzgHH+0WvQhQ2vl2TEMsnTukeYa
krz18Xxd1PGk5M0oG0RmTWPMhwKwJsBBLuuuYn95le61hUAn/sCRCOkYCt7893E3tXMGHcTtZGcx
vihw5bkNSuPpkKAVxG4xmIRwo631qSnl2ikpgK4FFOWhp/3fYTMeA/3YPiFVdtVqIhcndMZ3c3gs
Sr37WCr0U6/1xlUcB8jFZuuvOXtTBHLX2ctklm8GuP2N8XUtbGh+42IvanznjdwoVWNHWCBeePP+
wvm1Qpg91W+gv4BkPG9JThL/vZj2m203yxSNI6qkU8kw+aNbGiN97F0Xgj7ssr7HLDPbJjmVbJ5J
25w6phRgBaNxVMcaPcgrhezKP/wcQ6CMdLPNiSU4QdNKQz1LpsJba8PSAhzP36hZNjZ2EygZCUcB
XjT5tPbsqxQXepvGibi5q3bR3V/8TgJ4bb/N9zjgkCkuK1VczDtgwRZzj7gzNvZ/iF9jGfGC63av
QC29EEcjCAo4FH9JrVlYNVqbSQAIvPgjNup+TsxKUUOsysaxY5t36jS2aIa8ub10ZIATvlTH+jD3
TPOOXT8Ne+RY6oEro2XyQfuzK4O9X0ERtshf45sX8Bh8wNCL2x8rfkQOyNX5plh0XEzi1anXc2Vj
pHXz38ve1Iu1E1HUg+4gwJ/UshHfaTIu3l1kk+0ihVMXxIHRZbmQzd7H8jjdfYrhZ8Rvvy/uz4t5
UOUiWilqvEdZvt+XQ1xTQjS0I7O3L9OJpODWrlhDCoc6gk9q7dzI4aTmB9miq7QWDqZ9PqRa15BL
sUHHGl29GLia1L8AiUwxrCqGLSgwD8z4O2iZ5U2XyUNJOyKPrgGc0sud0h7dspTkklrDnz8MRnqC
hkSlm+tBuAL30klGpG6kd7mIEQ7+5KnGJTUxvhHQjwnnPbHEPVIeuHWJgsXfmB3Rpr8uyGeYju50
q9Nho/k+tzQgFXksfDfYdocKLAxLk9XHuHeieW2P9D0EjKzwQJgf9XZauZ3BnlAtOcc9G5AGdgLn
tpdQBFQRP3zsHhLKv79u6pOgM7LoVTdzAqITcitEWO/aqj1qHXflQQ5Zn9UOappv2FxqGDh0LPbl
+iZARhRdVGv/X8lz0X0/7DKhETjfN5OZuGz497sIsfJKBAzhiIlqEilbb9l7qYuNjrvuOjfl98SB
WJuTcfOXwB5RmWhHcxeCNvFG2SfDcYD9SK1KtaqwhWmL1kYH96b16s0rxIfKumZ3rGktvT1gUzb+
JdLhllZSfEVzAT46MBLTLwJ+Dzci63sXZEUMzNYVp+ViKH8eKfPfMeuX7AjulSkEXUZiWIX79zAl
kXzZ/9TZwgN2/mZGsZrPygbnFXa5UwVU8/jwzEtCqpNVxHySwyxU09PEGqWS/JjQYlerueW020QD
SYbLsu6u+01YwHpeSNR2+fOGtN+OCcYx0opz2oWTDepWah7lmsbLFvX0q3COpiweCziCl0lPcABk
arIH8J7kwY2iJWpmWQhf5nR+evjeCbo06ebMuA3ebRtSXYrCaNh4ZXR0cl9zFrfvdFuXgdcRDpre
KZOk8Q2eEhqcWOmcLF6Qvp/I+TMrkn5TOEa7NmexL8bhMz2Z1pzCxkd/Q1qpZKjcLkXqMFhE6MFs
bcNyLs+qGo32ycrA6cGaS4gEEdOuLg3+qlZRdQ+W022sSggKnlrrXD9JpnawtHZr1vH+vqNzqQ3O
u3OQQxo7AjGZ0FDYNWeci0nN+hi8++9OJo4XMoS2grEHnNPGcu+ZGoBKobe5IK0qHfdohSW/MgYI
GX2AlFSeWAtkwoKTTnBFzQEtHE2OFMBvXz5OBHhTTr+svK3DSdRNNWgzrCb6LC3wxDU9YfmQ/TfH
VlUgnI2I0uoF2/YjCL3pHe6vJ/XgWdZKNd4sja+fP8cNO+077qkF6el7uol8KEkk8Dbv0dC+YkrL
mdvS2+zKGxeYgrRUer9T7ystmxnu5sz/BS+rxdY3XQPUfUWHghJSghkFGghGPaw58ldrGQU4BxqJ
ikW7hWyMvyPl+8pvRSI8u1VUxhW6DGz/+z3kIlbTK6uSKscZsxtFu2fqA49E89upB/8CaORlfWvC
o0Tahr0MPQr7/F9vhFrGJgJSvZiPKbQrrLiOAkGXfWSzu+TfIbdppzaV7getiE3cFgKFNt8C2Rof
7ktmT4IEgW3HFKiZQlN/kWUXymSyDGWNwkd9euidEl2pff9D8MUJmbeSVPwHIvzMe71iyegdBfKl
R1dSpVwsmO7RM4kEAPerVaQHN3hqE/58SI/V8iSkE49/Tlp+3yO9pD0aBhYqVEnZ4H/GxG2mFFdR
fnlny+nYSIWIzp40vmq+aF7DEHxVYtnHDuY8N4Nw5GrsXYij1DiQPjVJw0lsR8az5DdNtlywttdv
0/5XktS7fLbIGR3EJcCSTn+vK14UJMZloSAZb1t/38tL4xo7Bh04KdQ4oLpFy+d8D1ywlOcEnFdM
d0NGjuW7K5GNzYv2+/wyvMRqT61kSASnepTkYDdbafRlFFIIVvPvj1uAlR4M11s8gGPgTvlEsX6U
FKi43Vpgd1QQ+vnUaOJQlD4kLSh/JjQVk2s3Ov5Z/mS8Ef42qEQ4+ZJyAtjTVeq7tmSiAb2neHEU
N0iu/TWAKEPPLEoGGUEP7c82XTkmTAZwzP2nx4fV43/camUoUuciC5aph7Mr8G0ZCTyZAMPto9YG
E+fG99jF/WgK+I3V1dKRM2PkNhfmXTk4zfHiDvC5nFcQ95uK/F45f1Mt3XNJOVE6UGRPKU/ayQR0
9YzKALKyoswjBqCCcJknxzjzKzUgnOtM/Z3ytj5yHuA2hI8Z0FHEu/gfEP5A1cQop7LOcebSi9IF
BEj/WhvGtt9J8jfufKSmHm3Dxr/BEM+Ud+W4tIJHnChctku7Owxwm18SVufDlxnsgp1SQ7+ghfhj
kHI/Lo/zeFTXaTTCBgDep1Ypg4gWxrXxt9ZBZv9vJTX/a5pYPprqQ+SJheEg0pvw7VhbEfd7uWfn
4wdK9/cfgnfUAwr/7iNupa/2bvWOPUKEYuU28gCOkXzCTdAN2Ntt7VLHrFWJ3v4yx0++TUUbJwZE
asIDdZhuZAwuyQ/K+yJaSKs7TQsnh941VUqfiYyRGABouzK6U0C4NYOqLpGVf2TnXw8f5wQEUuCM
THLpIYPLTu2xmszE9NODdKK2/hhJ81ogLAbov07cZTePEyoZwUeEkGyrpIPqPIjlikUFr2hChITM
5sC6OAZuGbrJcvbfVVEe3m1i+GbEEgkQ5B1Qg9tY2mRc2AYcUXnGlj2TWulJr71nksrHpHQJhSCZ
hi2D4bie07ftOAuiOxHgtmb7DAirdKJUGFE1/LIcrOLz76VeGMCxzH5J4ax8ocfKDbN5ndFYhnAw
1woWPydT78zTqyXluIjPTRK4LneoWjQ6+2qjZaG4BQ2m0JvRmLFHG6ki/TWyZ3vgIM7uSOYiJK2J
UmI+ten6Ffrng81CX+neyAyKO9nNpIqUNBoz8EQKB9YjJ7hH4rJPTV+u/g/tJFkiDcGxLA7bMime
XVR8qCOq4VWOC9zvejynbewc9Dgq1kAVJG1jY4EfKhD09zxhRR8H4TILJeosXm+RpE4QRtDxfmz9
ta0uZGGDPEbbOeWjSCNN9UXGMjlgB5FBg4Y33JV0iFrTJnxr08ohKUvydfwR2lnKFtcihIGhD/rw
9r5TzUlafgImPz0gB1tKrhfHFNXWg9wwRgcA9vuuLbF6LIZlxW8izNTaccA+lchWc/1Q3tdJPej1
PjaUYMtZgxkwgF2cTUYdRI6dc9jW2ETlnRp4GsOkl6gr/5epze/rWlAtis2YjabJVW7fRIJqyNUu
AWxIfg0e++1M6RdNOleJjl4DF2+qUcpR40G7xz5Oraxuprm4kYwTMwmFToA0PnS1Q2OW1AMPFYo2
kXXmtQ6C8jExYyBUjl1EKHYlpYMBRHRbnukIotE0jE76Zviz7A5oq08Rj5IT5V+AL86+nFuPaWV/
eMQ+Y9TpAIjyrYoJUune9HvuT/psTCYBzIYS00c1whDNXptqTvmcOQZ8BPIfd3nhAQZqPbaJKMcY
TlKsiArL8rcZtIOGdezoPlei7EvwjiffN6Mq/2IA0BTG1rqyWwj3K2c1O6/N6zlbfvi69dV7SSTq
qQhlotNRtE6yHrf0RPPSl/cHgo8MeTWCm3IQLCM5DOZ4nzgI4JRPY0l9cCx6Rc0kIb/0UuYLS0jk
wUu+BKU+HER0HV/oxWUt9PNI+3rfNC9zwIbGINDCfrNu/ZG9w1TqiVZcx71qFlNiG/snT5gwSVYD
Z+gmXjyrx3gymOhaHFLsEGIn5m0BAwD2YH0cUELkRXdMdLTggvF+I0t2VUub0a3jkiKUmzQ0qLem
wMJnK10kSjxuqtzRvEIRIZvsBKwDolbXTA+VbG6NHXPJg20n/3zA9Gwt8O1kpBvdWJTSyuw1kKi5
ZsC1VWW5CxwTiA0ryf38cIwlOEGF6UTX+QAmJW2CV1oaMwdn6uYl4hXq6d4IlDBVT/Q3LzIj8Woz
ueXh8O66W6nIHxFqxe/IPnq1xCq+ISJ8CbT6u9YZ43OrXlTiTPpJBhoSzvf2NMg1Na7veGamiajd
kpZSLFwhFsnfLsiWyeQRPK0NicLGHZMu8o1+MBim75PTWjrd7+BrIUpA2iLk4bFV7xKOvvW49+lC
3+vSais+hKSlePjDFG7BeqTA6y0qvG5bKtj62+3EYQ4A2bdTf4sbO/xLUImaxEkBb0xcKI/SnS20
MKJ2dKgLS2wyDa/U859VQ2BEIaZJEPdNU8pqesqQ3CwU5L2O44nXqXWpyoPfwyF6y3rEI+5hsqN/
uKVGj+HLy+sQgGraa5dvgyG1C4CNv5xd0/2iGlE0316A5MRfgsPe+f0h+w+ZqVjCeHoxCq4z7oe1
CElU19aAOD5RP1lcqGDHWjh1MhtOJUwaIIXZdYkBpis7nlZQW71YkfriUzRUDnrFaSDS2yKy4k/Y
rO60qyl/j12vDBAejD6f5xASNef25ntnqcttjKVOv2aMNarIRpStOaqSoWrKGRPjMuMz1WhqdxCi
rwj/iCL7/dQ90HSmMZRfpjY2mTcJ+N7mHUJme/1VVcgtynNvSzuPGLamOVkRj2YpWJg6elcDdmEg
GVFN2Zy4FJ4KaEmyoRGuENoOp4Cz0yjTD2OKfEqHBwEPZqknv6x9GIAuRqac7B1gCSNIAUEni6tr
19smT7ukcbBfxNI+ek5fFcGweeuLmZyX0O+x1PQo6/nfKVWKgeLTp95ScmOKzIOrMQCB5NR8/fsi
FWwwjY73vT13fO5FacPbYcWt1cKixWKfeHSr/9tRUzh2l+Zs0bg2VmFZi82F/r7bObEd+I1aKfQX
ks2WHzMAcYR5csj8JOaHsy+M5ImWYLmC6VEK4IhxeXxc/viRZuH+y5zhCjOvPDLeULiK+pVAU1fL
9QdC8WqOGu/WhTN3bA4wfmIIN7Cjf+hhejLgW7ly7FueLAjvqizbiw+1HQQYWgf/ZQ1jThVK3PTh
xTV3H58o8Dagj1SobK5H+PVIeecepC9Tsue6NNPsefnTjJQS7tRrknu+bhKkuGyYgApitH3gr+ee
jJc4lxIRu1Q97H5L89WP/72E2YkdA0UV8qiP2i5S+7a0LwVth6WdkUbEe5b60NGanx8r+qrG1IaT
W+rakHwcKwLxsi7SQVJE62y+JiiPiJ03eN4aexgdFW2DQlA7v5iwqlS9BwdQ06SMqwP/4O5HUMXv
llqMB4AeD5hIJZMwzNhQv4RIF0xBL8bjjkzPmNtJU5UiuR5rPURo/t3O2eC1SCAdvr1lXzMQi4NV
qhH/pgXKShRY5aM7Ut1GtWi9E/tSZzWMLwau6Zao45+AA26wTWe86gB4AEgLUZfzxZDS5NaR/xO9
pc9Ev9vjPcEqFEDK573BPuHXGryYxbNSKskrY+oadNVDeEpX6UMdKIumxvl/Hmm7BcGEB3R60wj/
KexDGJu9v0l8rpmIWZimhnbxkWHlyV9Asr6hNkefCdxzOjPqwktUzt8m1fIz66PVhCo0otONp0rN
27GhoinWMwCqvoL31F1ckV/X9vopYFgDvaxMGIipJy3ywjaq944XcruENq7RrVTMpKIz3CZO9hq8
czez7DLgTlro44fJwyh4w8RMgX5A897iuyUITL/rr+i3Saq12EuqqfRKjBJ3ERXbWuyv9yCWgp+e
Q4ViBSJVV3U3UkxnUUvf6ykF5EGg/2rOMPPROaRvOkrPRBQibwHgopW1DrCb9XlHWtDCgRjFhLhf
qhofCtQUWCR1ld4rsvANxWcLOUeaaggBUC0DtSZYNL9KcZqcBLHbi9K5KoAFouXFMS/ceX0k0lyQ
J4sqolM+C7ketKNBGCkGD9eKAVCalWk+Jar90z/n4oVuW+kf3cXNvI9DtL0qAO+VNFChQy6Qqb6/
wU/hhXMzDv2r2C+4D1FF793eDFla/NUKRPAIaJA85I5VXlkNnx+swUpPu2ltJAQNSyk7PA5HCLyq
c/8tWZ6MQi17e58DLnkt/FFIpng7uXKUnvIXtxtxdu4RxYUU68j4V+pgylBWzGxpactIklWrXGHY
bfHAqnqon093VaW6bQL0wCbrHjiRkv1PAAUY+hNDUEzQonXIaAxRKDpQ6JHVFqQ809JJGvAPvTim
zd6rs+BJWXqG1DxgdcesOfOsD2iIZTd6yvbJp7O44ZCExxMWLQdMQCTf0K4LnMF/Z1AaJWL0hu0P
lxKy7suFAZT5/k2QMPp39bMrb+e4t2SBckji6nBi9SOZE+kS1quI7WMmww0jDTd7wB48cSE/+/JM
oK8u2Yh+RWo+0DAOYxdDyGyntKiGzKY8a17yTfs3EBX40LwDT489AmmH5N9jko5KiNev5zYFUlmu
bBw8Fp9iH1he3sNQLG+vkwWTjnYwv3YGmsTHXej/EFzLqTcdy9iDFrjk/c5Z0hBTCWl+97R9O98r
2KPrbAdGPsDainq4oWtlgDsEfKl7P/m7deWyF3Hr958W1oBfbVSjm7vKSPq8ACrkfAOXQrMzJ3Xj
SzCReYNfHsd33ieFvSrvdG+DyoPC95KF2Ay9AhlS0H36a0g9K/iDl1NZRpNA8pYKU4ulqc9LUVwE
70n+PhSWqwXtafX3H4VFua7KPjeTJZVpOm6PSMFY6t8eadMFBkDctb8AT2dyJoZ7hFLo3SgWIIev
R/xRFGUPQF9mArP5iunwuBaSFUbQE/cdf0J11Xg2xiFsIKYPofdqM0NBTXpb+M2nwCKAYTQlHt+w
fIE7gaPfYXe+VdBwM0HlfkjrPQQZ2su1UXoXTXBcYtWGp1FsCizpjphT6c/obzqnUh/ezqgiXvcv
VhQ4bREE/ltlhNb7UTeEZQKdXVF9k40l69TyEY17njSVLP9j0lNETZMeQKiq667Wq9pRaSY3OXvq
LGeMWEEnSq4AzG4+pyZ74hR4aMzBFatVH9rUTDbre+5hHrdfkT9+XVH9U49lLfJqAqCwZ7f/81Pc
Vw/zCpvWfW7iI6AkW9C3Ua8JtIcCR8+Gol6MlNQmWFGDpgl6fMTzgyMP55yal1f0NSCVWYzrzx4x
aSKNT4Y2ILMVa1zyR5hrxEztT9xrMyhFIjI9WD5pt1MIa4XVE0wzXRQwFVKZCgZ8EUgdcyNnmm4a
GngYV2jvezCIaVX/07E0aFkZZGG3xWLCXo2AchyoI4oTbkUT7dbRZlidxN8/pBBSM1klaBJJv5MY
m6R7AxLeKop4DAG5YY4dVGMqmqfuJruz2kYBxW+FRSXDJADOEpleS42zgtRpePCQVwIMiXA9775C
3mvWgVjKwZ59aW1GprbKXQmsRItqmcpokqRJBtduXeuarCuUg6ESa+XAX5QHaffrMzsIyiT2ruJi
3a4KyneY3V2JeINXzkLyG3HOTfs7HiyXFL9IiKbtJJ5MeJe3F/fh/TvUKNYPT3DcetlIwZW4kc3X
7PMcB6Gbt1W8R8VdtKME0n3VXONTWYCiUs8IEKDFbwfnxxOOlF6iXZH3dSZYoAl/0hTN7vEPkOaH
zIfNr5vdjY4jva8rtYer3Uq3ezW7tqrZbIL9F4gh+7YYMeFs0qX3IVO+wkaRPU2fTs+KvTWqlBxJ
JS4/OsK3BLMHg8e3S4nr9VxgBPbhNy7/b5aLOpGPThZsbvPudLMWOLFyrTGuI8fvcyDnSxqVAryv
eHK78ENsXr7vV8Ir77lutZ0IDmvR3jN6RrJR+vpepyyEmOMOBQ7KfOOc+BkgdjET+Nhr4Shi5Pvw
cjrXtGW/OyOVuwZjOVHK2XgBZaqMIIDMe001VFAf01CUT1Pbp8l6gV1FJolps4nIdLWWK6IvWq0a
Dm/IES7rlnS/tB+rXJLjM6u/S2V0s9sDedFhy2E7DIYLItFS3KXmeaYg2znYzQ916aH9hekml1DV
bAReLMzSI+Rxq/8/Ca8hm5hbFsC7Q1sSR8S3Vgfxe8yfYQxKlUjI0YQnGiTWLEDtASbNzP/Qn1Ya
NGb53JpHlSzy2A/8xZU8FwrYmDtf/4zd2ab4aMusYac8RjUHyQcfQwLKgAaJ/frA1RjHBumnKqED
UHOX6IMOHJ2+LShsthoOt1tBJ0c/vo5gJZ5+B8tqq6yjMUg079qFKAJKF/BNQur/1KFEg9mpuQiR
X5vZiVsjeHzjxR4Ic+bozsJtu1gWvibKgMexYYKaKfeIpC9Wwj/cPWMAZfv7vdXUdt3o8H7LSyG8
cEA/KNDBjtlU/EhCIh8jO5HeWFodbtWyqvQ5ONQydhxlQx2h49eM9IPHQxx1kfGy/h5GWWgkUsMn
QTfYoAuYYSJOQ3l5NzXnuUyHn5sRwH++CE9JvJU6X9X2bf57asQMqaynLfb2XdKiaBFIocvr/zfH
VJ4quy/yq/BNGkKW0VgySo00eL3ETQsKp1t7Gi1fi6Vq6G/UgclxU8DLsTSWjZtUhAskC8cLbrZb
Ah7muu8vaSgkbTwupbGi0AN6qOWDXM91ZNc9p6kYcJm4l2NMSfdeWN2tbhXM4D+U9VU5ftF0/MWC
Rt/hLlHRrouhkVF8zH5gkVfM/VNtC09kMmEZg1y12Q0qlRc3fB8HGiMexfBMzbfQ3pMmF8FpXjI1
DyYyeUp+e7tqN/U1sm/tOlJoHCPOdmFrNO5fpXxobqRv/JpdibFaejHBEvtVGhFqUWf5wrqsNLRi
s1buUDD1sefKKUYwbyT6XA081sAIpt64wahFJ7w57ru2FL+0AXuSMjtVIHIGVIxEWOggBGi9e0w2
QD4wgIQziOt9+ZmAbaiWdKE13vMEeicSQjT/VU1reP5hTENu5Rl0WQBG9nv0AzQUcO6i+w3HrTIQ
gxBLLBBiquux01Skiq2PSaVn+/xX0HuCK9oeW0P0/Y7vOC5ym/LZMSCyQqY23/b1iPGeFWQQcq2I
g/3rY3nmTnEJHWU0G+HP4agjDXK7vLUvoULLgqRwQHL4x5tnk9RUgj6/eMM0U6+y/aiZ2bMXD/zC
GCegMiIhw57ont0BmNow7fO00jFGTKsw4x+scr9lh1WIY/mbmfUnR9Tcd2iheKQYMriPLPH3ZK5w
RYsYDSsrHZgMyADzG1ZTTMvS5G4msSV6YnPrhZfKxRbAm3R+oJN9U5os0NDBnOfyyBIbuFi8H6Lj
eAtdw69AruO8Q+VvAtuDhzXwT8xMWZMcoYkGu9sfU1m2bUsl+UG8lpQC6FhQWRueUgOcxmhNSJz+
bw2Fq6wWFNpIukWAdFzRdwwRMSdjzB1v8ZqrX9EvijSPZj7vGgBA2VRWiZ0zcGv5lHcpuq808nWP
T1o4P6BaCvciq39GFwYgo3yXVGR1sWx9CTkwsLpeWoBt5qFiE3H0+XOP7pU7usVvz/vFhB5v/48x
cYM1uLc2ckgvPGpSsHLvx0t8I3e03E+DIf/XX+MQ1pSpNOdqOE4KHRlIaMwDWSSL3SnnD4QlocxA
XtH6TadD/f1uJHHE9yvb0E61BAdB78Ui0+YZTIYb5+aVZPjZnJ+TrWqIscGLPT2i4+1XNa653dzH
b1oH+cm2U8e5yKQniY6Q8hm2/TMTmmkiA+RzjcCEHvXTTHV9cQHu25Jypg+wb1j6cKUGU5s0NZDz
W4shBo6gK2UygPAGhJJurJAxoiZUos8sJH7fcKMVtPuUjys8fewbhyGEDSxzJVRuadaq5JTmf9DJ
NFojKOWSUO6u+xBnFmyZHV/y89IniqBN5hdRzhU1/Rd3sPoaxfRO4MZ9V5hH3EHoaM4tlWZpPhb0
bmJxCD3/PebCjs6fMEWLlMVYht2hiz/1lTChDo1W0AsjD+UEZ+KXilisb1gGA1p5K0pMLMvERYiZ
hGCYLtQF7R/frasrrSTZrE+Q8vDjtpVFpe5AHtIFFP0CNjMHHAmqtMfaCsHTRWUDi0ZnF3efPZeG
EKYn8RAwD1Zs211T3hLuVjWvlWAf6y/mlelZuSPc/B4N13M5wPhnfsos2I8AYjWREbUnWcX6c+8b
9CHHFOagME21uIPuEKnNM8eVJ/cQyBh/b2Vqi0VRWKDYsyZurN5sBjXsinyzEQ6d66M8enKc0MSf
DBjeyEeTJwXo0cs+6BuJr0UsQ28fjkUacRVVwALUKUV0wfhxIpLTQAzPKBEHkEtAEcIfz/AoKltF
jKpe+O0svKbUk8wx2LwErUcwpitlEUiZAsu8VBUeeogsSVpWMTRYfji3dzufhubDHTfEn604NTOh
n5riIbb57TDzr+pj/QpXN8xMw6ny7Crmp1W37YgzbDegK96WEF/CR4stsKOZEce8+t8lmLV4CxgA
Zt87Qc70Y6mezkM70pRfCNb952P6Z7iLaCobvJiOV59zME42aka2A4eEzo8znwb+ZZdLAyYylfio
YuBTFZVLTRmSmJ+9cSQRweOGksV1tm9z73P2xMtLlBD3tqQH0nVp+ydK0f+/GtPRO/0m8X7wzMta
ihBXDE2TqM4j8EnX496N75dyhYnry4awZYHekQD1rLn7if2OI1DDPWEtCKj5XfWM7Lx2RvzBJQxA
OS9MF4YEKSW+lrFwAtKv+Y/WeOISDA6s2SFiH6cxo7TKzNUEAmft6OGVr/kITZ0bziv3btiJTv29
E5t7UUS/Gg2IqHFHvn+pPdrB2zTkZF/xKyYNrAH5s/wf+NuJVTo5k59dACe2WQUW6XeQ9uDSugwl
qzDFukCf0uOZN0zkiHtIAFTNBn05mAH2ATTXuJIHmvvAGDu/jso/I/IA+sIECu7/oTYIbfnxA5GQ
g0URTdd7lVfNV3LE/q/biOL+0MmBmTfu+xKP49qlzA26dsrnIvilGFuSUbKDUB5PBdtmvzzjIJP+
V70/sT8GBeEdK6Q2XQ8AeDX7nf9LY9hnh2hRqfNEN5bCKAk2JZSweTXkICZnDwlUHJ8LERBAblsM
fe88aLZ4rZ7XDqQUSjrBArZdAyXLkfLCom2KE0adQ5O8y+Oi003mTuZKWP/Cx+dkqEjqibgOZg+V
C4nLLe5zlk62MfuIvcwO62YnYTifpqKy8WOWOCz4dhTzdX++Dny3V9c/p957eSaziDLDS6nDysK/
Jh3eAH9yeDBLNPNposekoO2tBiJwRkzOXuWMRwxWEDYW03ezwfwQkPB6WrJsmytcKmtvQACN/J1+
lVQ7fqzUrwcMISJdbXEXHia6ZJd0q6OeprKbyvCQDMuSSfLmZClBY15S2p+hodvPWCSPb+ObpK/j
tLVQTNDj4cFrtD1qFtJzX8OD0zW7wtnlFAPTfs6kD3n9oXbph2O4uBWKDrEOwFlt8yOfCy4G0FBb
BOEGRldMVDr5guua53xkep//0cMXKvpVypVBhjaxP1zUyniDoCT7sElpu1FbpVeGkQ5DT2oGLp8s
yBL4+WH0m2CceFifUxmxKsZ+Bonhg46NtzFmBdlV+NHIfp0s0ABEpHwU2hRkAk/rt4AcBW8HiEO5
g+0RlniGa+tirqOXcmSCAbp8pkKSPYaqVbDD+zcJKnkY0AJ8pR1fa/I32Rj8r8V2jF7pwCuPQge4
8L9rxqTrLrD7Zodut6+OAzyG/AI9xfQ7Cvh31EzZQ1QJV+vU4NF+9yrVyPw8CBC9Axhz54fGBjEh
kfNQpiIGezWSDy0xzDe4iBSzlgdTnB4+eAKL1+dBOE7to/eMza+uDe0Gdo2KozUtwIPVPOATuyaa
EtBe1iGV70K7Zf22YcmQXG5iyvYI/cf2QMyQKCrnCS4VbuqXxJ07OQVLFZIZS5vbucYQic9mhMGp
gwWNGx9wJ9cHUUmZlFDz2oj8Qo/+d1PFQ34al4mbBWILSC19DWjkq8RsizlFAkB/TSS2TpcBNjXq
c/9HaW/9rAapzFPNpRlrHo+JaI2OmNMAGv4qrMiTXowhZAePUgAiKQUCsjdwZqJ7GeB20YmOGggt
IN6CNbjLJEr40I5/rmG0/Jo/uoroBvYFSMAaGvfvs5iorfBz8eagk4Pe39P5sSleV8ky6+eOfu+Z
kVWPtACg2PzXANAB+QehVMd0twx5b/9Qwe6WP7EyaoHeQY93YCYAccSOJZb2cYhgOJo0D3Lv50xQ
H8Rpc81lZeMHHWncRjbBKi5Nu3H977WHZD2kitVIU7pOWMadNmlPK2stt+kCmzOayzIeZ1eQEcq/
6CocRxHLBAS43Hnk2YihTwKqOulJEBkjgvn3EIQvvSW0tUHav+K5cIb7g/3HsMV11Q4kKtHrnYgW
LFtu8hFmIxd0Qm89dM15sFpFmjrfRrmL+9HIG+C62oJi38itvIjGrEhZrQrMJlgN+iitowIzO4NZ
fvKCWJNolgtL8jvAxblHmSjievaUb81Dqd8+9NpvXu6i5OIVIq3GZvLgwHPMOFiiXgDGNySEdGxg
7smQwbdsaGUTNVb2OBR+77EaauBSg29+/LzpXSHG7a5C8twC+JN2BPb2cLFMUn4dKyrNXXV3iSIP
pDy5UdqegrM7gjehBO2r720MmoNKqpnnNoYnENH1f0xQUZynypWwxmpOBJn8B81x+VuNdtuL5POj
fT6TEoYJa7XlsjXFJQFXxtgqtgX7LRsGM6tF7lYmoMLjtuBiKvugmbcn0GGmrb0V/0Vkn7Fp97NR
3TGt0EwZuIZPdcs3UFZYJMUWAl867BDnw6xqKDmaIAOfN/iXLaV0SK8C9w7xxy0GYBj5W71vUUMU
tYfwPmZLrtNtMRdePJHJHIxtXL7Wjtx9yvKU8YmMBayh4jRBEU1s9ueNLo7++Gek4WdP22h5mcrA
Z2dqGc47oBXt9S9LqfqxfHYa1CAgX27ZzBG7oaHNDFjPNjrjfWPvC/N68E9iELBkjlbHUXsoKeMC
0M46Ohj+qAo3IFGnK9t8bFtK7RY/JsKSf/CP3RmTj+6UpmYqjaWEqCat5BZnJ44XdCjs3WDjZ3ra
l+9ewSWIxADPZBONYmhawEWaITn09Mr+WffW7KjEE5zYV2x3csK5Qeh5TcZgeKpFbTU43b/P7Drb
zLuKAqjm/VOJ2GJZvBoGYuTj36zdY1pvSPvYWgKvuEalg99F/6kVekSy+gt1TSstdZXDMPNu0sMK
pC42NvMSq9VyImlLZlM+hK6g/iSC49yRxaaHe+IgoCu8K1LXOO2ApSL9nticqqplB4H0Yge+9yyJ
WsMJAA/t+ZeCgae73LTl7n6FZ3DeGUSLr3+3RUWXjqIKjE5m03wONhqMfgWdxUThIuEL+aT9rWXN
dAi8DcLA8NBd2xiQlzQt6Sp0UyVwCrOUeshLvBGhfv+un1sBw3BE/sY12AvOm0Ajbfp3sHWJd0qa
OCvDGZWYup6xh2NgjinKnVQ5+sgzWSiKZLSLEse/lqsxQCRcph9WRTGNvDybxJ3h+vDpu58C/lQr
DefarPqYblIpoRX0UQ1y7hXXXV7qpOBk4QL9D170q1Zb9EStnJjhAxrn/Boce+WUwmeK+TjNfjz3
/QzvG8DqEUyExh3FjVFq0ccCpvPlCpXbvu55j3IvYvlSaL49YY9FDPd7QIRgexrTkwCoLnowJrhP
OJn7yNkGpj+XdIGjZ0ZP8uor1R8i2IdjIlWx9SS+l32yKNEkq7CfKUSKuhVYVYdQE6h5892CdQ5T
fDgp3NKX6etGZ6wqCf1n3T+VbPYdDGcy7PIXKTwh6RFJ8j3ToFb40sCRnHwR9hCvj1xSnHlq1ZTe
VvDDJ7PgMclyoN4RxAtzIwiby7c9Ub9aJxZOdyOmbrtM6428EA/6qwBy+/AlHX6kBYwc4kG5+nbk
c+4Jv26XZE77nGiSZIOkvhdhfhwvMBH2KsY5ljxHtayfQIxD0V8UWJNVik24gKxHNAlHoHux5FnW
UIVpQfcwSHA2Ktxl9F0sWGfxpSgrJzr5HwTSbgcBRK9Vd3jire8pQ5KYXfhvWEOvf6MrX+QdQq9w
Mpjyyket3Lj1oo8MHOOlMt58HUn3JquhH3cjWT5vmU9R0kTk2fqnblwRwQ6SU4rvrHH6sSp5q9TG
yFnNR88KEF9cQOSfkt/IOY4Mpx2ez/s7ZcsimOhqdrP4oeXul3ZUeu3lrCQlbRI+ZgxI2pDL4EWl
peQKz8z5au9gJ3s/enR6spNBldk8HqnYO0aizfTQOSKt3LsZmE6zzshkJfykCzkFZj4RStSAcxny
xNE6DlBclzcoBNI4gATb14PnTjEtZ6R3+S06uXS7cxDLyTkmHWFCGxFJJuDI/iX/+lx0u0F2oXVy
yy3ml8703ab0Gl5WhkdHyOYkCucdGfrwOFLSSq43rvHoEfvpycrXPCb037siq08MF9u30KAG+NTW
v5NZb3A2YvBN4NK3AyITmfs7uoIAd5/ci3/VaKKpDNV4x0JpZCpT441mWiq3uFtUKDmGztSh19Rc
EIW2QRjcowRa3h/W09JuzTjjX0TzW2iwSpPMpBqm1Xh/u8+1/Bzx+Tl/GLhbwPd1QuSWhqm6+Ews
HD6xIAS+aIF9xmEpvcdYB1CwjFS+ry8OzGEjsWNdMRZIk46WVDg3xoP2cjYzBEGrHyL0VfqbLqNk
bB3dQmnwAw/3np7kaKrItxqofI4y3v77vVOgrL5ABssdxAC4xOigbLP3QjuMZksIIYaNUi7aEJ+j
3P2GRjna0HkRM+1YtKA2GqqmMygWcgGMr+N8NRoX7XIlgfcS3FQDCWL45NbWqpL882kc7WzflMlJ
VghVz8zDqLMtsILDuGwNADCmqiexpnTZ9Pl7HCoeuOfE0LbPSz1WdqEVYERSz3uGttxDdh4lxV6W
m+KmuWa+vWOsSVK3Z/ARiEJY0fLMeL+upSSBVbExpT0NuHD5FLf/P0NTTDHg6o0QB95nend8fek5
gngZtWgkjoFsrbUoPXCFNGlmDzxAtJSVaEp+xVwPTCn5lWFO9zEG6p3zTG3npivdZ/fACPMa/Nid
fh1jD27FOwHkkGIUYO3PvYIJa+Thjfpr4r2s33u63hzN0QOPMgYsxuw39IXbpXExn6x+QUd4YNMA
lWtvOrIZBpcry47Gc3GmoWAdw1BUcWf6zOli0UpbVtG7YkfbQvNYsWzMtFvel94sixOmRrniGUMY
zaAWAyXOVWJ+qvzYFcgZ6mP7veSBCLW8q6azc+9rxDv/Qe4y59QyisWVSftFnboaICo7mpEu8Ud3
7Evt8Q7jYf3P5gOP0eYUhRSa0uDCcXR2GcQiak54njeSPt+31xC94c2z9iY+z6rpfPmijhkFlsUY
g8vZGfvu9MjiS/KCWRSpIELqc34l1mY08rHKQLsKYUEOvR4LuEJrU6BdDyxXNF5YvCc/V/85y/HZ
EIy0EHJ+bm1AUeHVCyL7UIPpcLaN26WmzZbasAQDWL/7OT7A8M2nfjU68kOVxYWmOoieiS4YcOpH
fjCCsIkRXg5otAPKn+ofNM0+RX8QY+f5BPtzJEuiss3t9Kpz6y0r0sfyzAdnlVwyVjC3q3fVJH2c
ExeWFd6scgsmdn6Y0aC49Jg9qdSKYAum0M1AWDCrdRYBHcDWBPrqSqwJxfXAj0alqvrAZiQyCVAy
a9g7ZAM0qHnnJjhSTL/SgUKUOGr7qVsu+A89cewogMGzdbFgmBwhbQAiV5KAw9IphjNY3nG8PSxq
As3bYMeXlI8nCUCeZj3kKB0qK3nHZe0EI4LXL1n6wJNW4gBpmMwDqKshOC7sf4A3gwGbjwtoZ/01
kmmdOmyuUZTdZql41uuW44ZISMuUeJRQmYDnFxSmM+IbGOPqg7hzoxYE7bcotVDYgskDr+3Ul1hr
Mv5zRX7ST0EmkTkDqz1yB3VTuqMnPi7jnt/HBvSlzgOA9o2Sc2Y1fVLFSUMWLJ8ahK6y3s54wj/A
JiLFUqZ0kz0Hjxiko32asOmWyKWQv3fBipDqfzGjskRSjX/Xkr5ZHlom6fV62vCs/4dR2txnF+QG
uUGvJ4jYl8mKGk28qRD0PJEbGTCT4+huGoAfPEueh8MaGrpTift1nXh+xqyVlW3thdaPzFASRb04
gPvIc93vPlqMr5ayZE3k6YlUKVhHrlRfmaYT0IpgMyDwnHCPLSDEX9JiAmqOIvjgBJd3Ljw8zxOD
NcKwlLHnaO0F45oX/XzhqXQOac6Q07U9OPPFOQxKC8IAKRXSaRc1O1mtIyTUjuDH4cpHUvzUea04
oDpFy7SJ2WhNYsRAAvJtEU0f3VJht2XwKZWuL3YlB4WxWt/wn9jjE7LIELI0HHb9bQqRwZvTB9K1
/+kgoT/SeBuhQTrjWwzj2/BO2sG8NWXmtsUwzPWH/FXBoqD0M0XR3M/W0E/ftyjfwoEuZy6ImFTH
wGcmFIK5gkdX1oIf6QxoHkXVqQ1JI0Vi3FwLonv3RBkhf8S6OLEG7/KfMIHikux19K5Jpvzi9TGi
zUBOfliWs8kxpMoer/yhtrTML4pSDIw8RAKctT8/dR+1FBk8NIhezhKoBhG31vJtpo3FxjDJT524
Y8VrH6xEXzAkolmtrpCzZLJxNbmXhSQcQLGy2t0K2vWDnpsuM88h38BoF8YrGFY/Yi2j8g6w42el
ZOLahYzIij3V7Xn4n5gvANfn0Ex8d9v+BthGqu2yOU5axL0In8TrGIxF48t2Cc1miKS5X0c33Qfu
9AVNEgd4DoVYuddQvyxNUviTiVDngTCCm7ti3mlmDCA1bKB574wjw/Km7mm3dusrg4zAao8VQhR/
bjOXEh5d0oQMJh6lMA+B3ZaRybFQXiEdR+JBXzvixlCVnQKyU79bjrCW48v22YPguG0c0unEfifK
5p+0t2EuocFR0JaMpbv1CxsBA/huQZ+A/wo9LKCykNb06IEWTh11xMvNFzNU855QnVxMnSIHiLwq
6l/aUJoI82B4mQN8iB0k6W50Ni8yC79Ls2GERKzP5kGuoF/XqPPinK47Ud9kBDRtibK5R/Kv7BQ5
KvgV6yTQdf8eWbw5h6cDRyOMaYLF2VDmN4rPQJPyfNh6GSo1zouKVRbEMmMF1jbuRMw+GAuhdptE
PgVwAtswgdJ1NyNaoAMQKb/PS1iPuur+L4qsvr5buSyiRh+0wVhh4jmHnNS7NFpbesht3G5xX926
tAXuqrHaYjUDJamoC6vfnqecIKYWEjKBESy03y3uc/P4eN5fwTi6F4jkC9s/xrXvaNL3ldlfa0m7
SQtEh+0Y3612DkJ+JzZhvDHjGall4B9Z0rdw1Kv4QR7fLNasP4Q15qpO3n7sQvB4lMzw52Hz+Oyh
Mum0J67g5IvWn7HusEJN7LuvK3OY8YoWSxgEJAXE9hmmxQhnujKvMW5xHBaVWmUzywKcT6ETKibN
mTooOfsbM4+wGyzTUYonhT8jJnkEWaliYpj8qlGzTIc2I6LX3lTk9gHGHrOGQ3kFWW0rHNSwWFZ+
5kPCr1hvvBbAKKhuWW0BUjl1/JMlD2dXGmZ6DBe4CssY2rbU0Ae5PKARtW6Aqm3f5ylmKF+7qpUK
oufue+0zvn40RBK+GZdwauPq7vLxi1m4Cny4n1JbRIBHkIA/URwxKEZt/fkEfuhmQ7tIDC/Ec4Om
T3w3xUzO+gPNlkb81BRpETIXKe8FDjg32IGwgAaUwOpoKOrSuzP6xXwYfmQocMSnk5279hWDyWan
eoKGSlfWxDv5R5+3APKk+2UuMr8C7OfiCsGTktrvJ1ykYoE/6owwoz2GvxxgswKeee8cszP7dD/R
WKjf5R0K79TgF1LZmtCVMcDDDcNIlkwl/+Jll50lIsnLKIfAO6ZEfVPKs2lrceb65e4+8E7MT2YP
cqfJAXtXuAObv0d1+v1vr/qOFCUnYW1OqgT7ugHNkS4k9m+UvMp9GzD4LCnwbndRY7oWIbS2uQRI
2upIAGcXfyrGUhhfkIi9V7woyl6ubki7AqXTz/zLuDRgUgcKChvlrRCg2t6hsNAE/L78JMFKgYX+
AG0NoG1SR3Hj9txfA8/6jDxHcCuSeFeSdkBq3CBLThjU4aDPQdgzaOvFB1PKJEV8YLG5UhKr97aw
A5BWZRQNc+i2ISSEItdAqnPhtI6grkDRO1K5xTTHLNWxTzp9z1FM4nztJlT/6EXmpjpR0ztkAl8R
dUQKQSjPzblXUFh1qq1XzgowFKRr9RsNJmgGFydaG6SR+LTuKgkqhjXKaj74EuCPpYA++8XxE7MG
jWp6Ly2mN0iXSBjQeag+H0kvpmCBhQfqMrhsxHYctFGwiQEueGAzauG4CC7qT7FKzHxz2HRCOA2j
wXEjlj2XG/87yTSLgw6R/uVsP6EyCG3nMjGVeSVSH2CH7SyJTWkQ4nUt9js8pvM6EUvhACLJpEAe
H0L3BufdJSpLlNTGdwNfnLlc6DZa8/ENmZKv0mgMAXQIOfvvXGIGgSDoPnFe8cFNytX9/TAdwRyJ
XlSWHA4+RgkfpCVRmdQRN6WZ3Mw82lnJI40LGaxGl/tBSRGzIHlff4Y6F4bL03o9kCjARoRU2n93
qGjbx4ew75dHRfnM6XtLKkv71gSAZAeoxoxytcxVUX8mjN7/BsSESYSdw0evRvoztp/AnSQpKFVX
hakWX3X3Ghpec44uEfr4GlFpO6HL+ZvczXxJwwmJy/LYV1sdJw6fB9+Vjbnnj/qfA0JduX1FzMv/
IWQ4YdmHwHDZUYQu82+xzwefdXSeBVE5qU07HRa/Mt+35rahrTyjfwp7cIHfy6KrSO8IlwhEiD+K
QlyXbguQDMdWei7ydSLzrYNra5y7yzKSLpJ20Hl6WIh3k5yI87LryD01lP2kIXeOmPExEr/C+Fp+
Wx0F5TYEGU2oGs6o/7FXV1PLVg0kbPkvgtLsVmD3F6ZsDT0CAWi0NkKDDN44zkrRIW/cnW5R0Vdi
3p+ahTH5tfd2QROoagvlcUz8c650pTEa5pl7vc2WeywPTrNlT/44zPqzygO8L6JU0hr0D4fInD11
Fc5vavngcW1TEVgDdfLwomYGMRLW7iCI38NfARYHxwb93Qu/XDSfpDLnnZPxpRt9FImDcpVi6DP9
JbFuIfGjR+z0JBnd04i8l1FYq1BNQS4r86xNlsUEsdR6VDn4KYXpmYujwlbtW5xi8e02qYHScrTE
G7+QjWky3juck2zPmt1XG8l8LXuiyoZ+Ft4HjkhqF/4mRbgxh7WwWnzazdy25Sk5RSP0NsEmI+5n
vs3+Xuuo04s/7PeGhN8MoxRPlqB1k7myjotcBgQ4nQk8Ex0EyVgyFblaDo8vTPWVTv8iUEQvsjmA
oqO8g+65MCgPVAqwB0We+dWIm73y585c57r1b9G2ydDpLBXPCkgAue+eH7vc5spjbIOMsiqfLbfG
PBHPCrg64ja9V6Drw+ioKlEoT2na2jqedSAR0pYzu9SGsJprDPwsn47QqU6jJ/6ecuGXQ2yGGoZa
+ICldfyFhm8BCmxN8udLXmyQse8Yx/QsKaVq2yw9W0lRQtpSNMSx9AuBI3wx5EbmoPSlbA+8/2L1
F5OYCpU6Gb4zWXzhSGmnSwkEsulvVVelpi23NmG2PAD3l4jCS2Cm08vyEWUYFGfHucm3QpjN9Vzt
uk507glrcJFzeNlEVeQFsll51pHs7qO1KIE9g6tP/qxUmtQPwJQKjcg1GXNfOe3F4lB8EAcX16ov
dyV89cWc2ZOYqpo8g/Qa7wFjnrEXbRtPy/+f8uZ9vboIOkwIGBnHCuZoW2wf17qk748GnpdkklWj
CDJ9jsoDggg6pCbMaPH3xkv323POoed8F6LnYNGgTZAimtHV34cweWvHo9mPXFV8Gkl8HOQ7hNf6
XAaJOlMXGCqTgP9avhylFpLR10nKhfa/k+NRJkTiAZMPeg7WGnmTJVuF94C9Q9c5lX40LpXdkZie
OBTEojtiK4aN5TM1Bc/S/5hLvn/vVFVe+j8Yw7lyyK1uv1cM9sW/8UXbb9ufdvGi5SkMldJUr1XX
TXYm/UK+znHirwkjJyNDWRebyVA5YW0YXVB1xrHth31GWCXhpXeMl1qoqVQc0fEe1tv4rLePVuIA
3gXCXCTQVceteg5OKd+2mbtXyn2hOmUtLflAovTf8ukLrkLwO5XGvpQSTWmiuY5nJVuzZpYxbpqp
SzGu5xkBlf1Tchr+w+LR/l3MeWy46oCnXtTGEvAx+A/kbYIlRSX2jo/Zf4bfj/DOjFZ7kr7E9tEY
LqOFjHt58zYX7q/WzP9vKL7iPiY5R+W6MxjlPGUSs5ZXDVEELcRGD0j+oKE3t2Xx5v11fSZv5qn2
BAub4rcDYvlPQFOFov6Q/UbdgKEaHkc7qJ6hvrUD6K+EhFvh2/OEq5APa0HAPviUWR4eOXRikNxP
g4vH+L1YhMmXEm6ZudRo+JPwKJUeHKbKWS/RAHc+lnBg6VcdSy05iWBke7ibDcu7GVr4Dwd9k7em
SIa1A5vV1ou5v/QMFn4NDpFrPw2pSRnx1w34Y7XQT9uXoYchhiPlo5AnwSPVsICp0mGDl5nRmvh7
6BNGoCOBZAVynNz6zZkiCzJDSqSSJVE8kxAlam4bJckuBfsYo+eLRChnppZIccKAWF1mw4iIkE/S
+vmWiKDlyG2Sb4cFXo3k193Fa4/rsSZEIaQ4bjVOFT56ZLlLF49/4X0SY2BW6aD868raP0OMrP7d
vBEmC64G+SgMKYqBBOEE5WULCHRp2jStpaPTZTxizBjqRQuHI9HEHGSDCnrLjqN46os3rWwXkcna
A9VwsLRJjUlGi5hNDUjtCXujoRBjR21v8zwkeafNhxV57im6cvlaGom+to8C9GTziYGF4NjYE4qr
OqfJZh9U5yXS67hCt+P8IRopXed4gfU8Mpq3ER2NwazcEnqj96Qjv1N2wQaPhRpeXoS7jHt6Q4cz
iacosb2UutGuB7ZlKpmx3x6Pj0SdTRJ3RUZG1tA5l8HNbnAw/De2BS7zwXMjYqZTWa0j7/YhCHxF
G3/1xOHMV7Qb7OH+MosBGH+Ofrso8Tt70VaKgZwf+EAAQOGIQaT812KHMa1FpBUDVbLCKBu1iVxN
bqJ3uiiMvAoK2joKndLAZeiLMY15xJ7s5m2n2tfCquDT+yiplw3TWiyDKKgePnjyQYZ2FGqHW1aP
K37/YJ4aZUO83GnLDWF0XYNOgeYymvLywcp9sBbJmJ4YrCeM3YVxMoqpDWQ9mp3QPqLLkr5vhhOX
h10+AO/kWR+5znMY/wYowfi3snUGTmUg8XzgtRNjKPedAj5ajQG7NkNqSLGxHo1wr12oKKGWHMS+
ALa/W4il7xD2ys+rhEmiashfk46R2OFRTe9ri6MTKp6Icquj86iNw/t17+sLk/9+Yb4Ske8xznfS
YtilgAZEGVf6mzWzS9mFQhRg3mcbdsXi4a7MiPQPZ5G8GbijWCJ0RPRrPvf0nD1uIvlEo0DdWZ8d
fSnOCz1V11elHF56KVMllBpt6flL7rAYUYmjnKizOns2ENLo1exCEeTRfrrS6PtSbOeJV179eHtF
rUaxAgQ/27ShbcJ+M7A4OXgjnlLuwCkTh3vL8x48i7waf7+BS0Can9GoWYWEXELQ2876oJ0TbHzn
006GvrYrXV69/viiim7R/Jm+c3dS3dkbzoB2TOesn3E/57ZSweeQbSvZZPMIEZXtaqkjGfTokARB
LhIr+qQ+Egg7GRA3lPt5zq6gplUb4rC/VJjZlIaHHB+r0vug8g/ThoEunRAKChaclXaKkqOw6ACa
FwLq4y61oYsWsUZd3JmrnDWUf5nSdxLmikPzAHlJqNs9pTAyiKkE6urtXTfHYp3iBhAyUs/QS+sc
ojcZYpLMaYEtcQAul/SHb2IcdkUJpdYvnFZhVPKAkNID3VFaO4X3twlfta7RvBvV/450poBMt3Uk
9kxkM2950JsKlTDQQX8JsKFd/Byi8XNnXLTCLGYZ8FZUHL+6H3nyY9V2+owyGwIfJadkvxe41ndw
0tA/rPEugYcW8SxjkB/o5YWtdxuwiLtdoJQCGNjY+eat/8Q4PUJQrqhykdB2OW4S6XeHhd5hJZUc
1FhHCwDMaxpHMtzN9uthVr9YcbwNtLCZOT+qs4wLGf87Lr0rtMa7JYaYQWIZsatzN4yrC+f7C85m
kuHJssY3s/6vE3ksNKcyu5RYBWCwjqNBTA2ew+c4MChXJ36skgjW1Sy7t79BgFtCZCI0xHlsxEYF
aOGVdwuC6NgEn3M79vMj2oPa1SRFf4Ru5cWfyjYpVAX5h6sZ1yv72ogN8FVRJ7g6IDtZ8kpswlsS
MmtulnrJE0RUvn74tmHmgE6gzDgBR5qey/vQWZXB/GLAz+1y3eMtO3JAPviEPlPLRy+twD0wHopc
BydQI2fnL9jScw0pY/It+soorHI2Z6mzJG+ddA9OI05kJbGY2T5Lo+TL+cnJMwaAxhTxELmejq/T
fVFEpxJp3te2yJVcQm/HZZkQzxKwtEHPR9Vl/tysE9I72Q6OFxtRrGB8cqlRwIy+9OFCA+UQ0MQP
BRqn6NFdlhs44uJEaPIUs+b0qB60gXR2a6vRQ5gVtWy4ME2UCwaQkvxcc8CbVW07OaSAhiZxMHjH
rIra0tWC5KoWQHSmeZvSvjNBSCJMHUNXzU06ZKNWozeEgpW1ej2g449fX3vw7M3Si7Gkpr9ASKON
v8+3yPRlii0MZv4f+DQJQOLDqn6aNIqQq8H3stVVfoOMB78ptHZ9Pv1Qa8C0xPce9B6VeWKb6wHK
mm1hqF7UNAZY8IVEDKW7eMIp4K1E6bPpjRuHD9zedU8t1lFw9Di4XAnVdGuWUGLZiNtrO68c7LRM
r+lRDS279X/ZWV34TuefC22LBLybAFMdZ/v+ODdoulmDuJjPECr9Um+sar0LfafaQaDyZyo91/Wx
dvC4MD9oUugjccoygShyaecu4qQHHBqH5a6vxNSRFrNBGYaYzkCuFADyOD2saxIDNPLWMVdDoVNH
eQyOezwiZx6wBNsTQ2Xk9MFsWSR/tojU/vK1aoUy10j6SnkG5uOlz8OmfcubTp34m9iydNeg7ayj
BNh7SjfW2eCoG52tMio8l688aCnRr23tJoPButc/sztGQQLNZliwYkjnxsF2dr189NFg2xO3ICFe
RKfKGmpH4doDlrdvar4YNvlQBwRU5YbmCKbr8ZvVBfhq47WCVsvbf01aodPZRiWzWhf6+sp02W1L
LbqEqs5ZGdrQY0Rwd+L5vE90MstJ1PNNOQYpFQflFA9Dhyl9iBZLib+62NEf1uMZFpsAjqnvxLrt
Wg0i8LS3gF1cjwSKgIJ5KNlusovrsjdsiAoHVOfnbowK3tw3qWp0wl2D9tSwONT06nfuIdW+xCES
xJ0BrURrCatQfFfMBdy/i1gQgh2uzn4eAs9uMt7pEnJDFyeZA+X4beR4yCTxxyFouTzhHrZbTkIC
cvSrctH5hxnnpe52/Mb/ssPeq0HHOM52Jug6f7o0qsuTbBOi3pVIc7BFcNkNQSKmtbaY70DQGIF7
a8JtlMy1rS591Jt5rKTIUOI1rQ2i6IW6W4bDrkndPqmcz/Zjpke7clkyq3NPT5EeQWNJQelcHV5O
loVNrTM1fyhoVGYtWfpXkj8TDPhN9SjnkLBCAe0j14FfoamYPef6O8p5qSLphhMkVXzVsy4e7vGE
1cuvCAkDaUrHNMB4JBD0JC0ItB8Cr3KLiya+7FC44K6Zj1CVh+aDNrj5JwnoxUn5ka7PWG0tbP0j
+lIbMCASAiuB21bQe+63uoZUgKx7st+5//QOlPC5xmr7sr411bI6hGlRS3Pu/X/XJ486dz/6Hnb1
shx/KkPJ8rRAQ8Arp2RRJWCC3mJb8vnGCqMAPnpAayo+lUOHvpjomRgjmA6GRfBfDvpz2NzUCFXp
NXQ/YCXPdvdegWdLQQehtlkiAZxRAa+qvb+RghMPEHpGohqKKXEo0Xr4byxH2LvrKRyOriOKnhJN
VhkZ9ONEuKowmdTwLp2a/wslZdYrKiRsk4tpsT1Lxslv6rIfVcXwAsoNuWU0JNZxIlxc7P87+nrr
+dzZuFOiOFUTND7uIIgcI/pdO+f/J9ipPte4eAXv0JY0ioWfg2yEN7vZMj6jQJjxA5C/VfcBN8ih
idIXdQHJRWeMbx6JBBXlyXqtHddygWRV0K4Ymu9ZCd6YRlS/bbUTnl0diDVi9o2vUpQXip7z9Drh
7GLN7VCRJLgHWkqsTd1QV32YbjhxpJqL/XzCCEEoB0UbNQLrrKFa8lDSNZom8THMpgYjxxsDSAlp
EnkUmU5viwVsoxSLdNeRCdsmI/1J3QM0VbLF0kNjyaVoUhBYkVPr0dPOUdz8hBay+DxonlcxOpWG
DJfpG7wxUdku/sn3kr/mWoIHqF3/Endyz3Fe7l2JdN6uId9fNjDHC59WegGqre8WmGWUcs6pguwF
bdqBWNt04RJcsAA/g+X1m8DMQ0xg8d+WG7Rt9WYl+LfPQClLe01zcX5kKGHCqq+zIOMVZ3vS+aVy
KyCRookTvpNmhEUHoVBGtaNHJmOoo3v3Ur2JsfnVhtlyzNbfSHCkufDX2cyTUsviE8VYKx2mDnge
/nGsolIYQUCd9HUjUSntEnxZ1soWRWWJKJJqJ+jI4+/Q7hwaK/Mc0Ns4c0ffCG8iKbLDZlBbhkLD
bpVE1xr47GfVezpJXhJA5LTGxkoSo78p3nuNbYcOLWEnhubKiT7FUF8YtqhTcEzYOFYscgAsJlSt
kpvZcaR7EspAl2k6LbIhTtWoJ1KhlxQ9YFeyuD2dBf1LGZxbKy33QU0y9RDxdMtciQE0LImn1VPn
lDfu3L4k1fkFYQe1lhQmaYPmxCGJgsa+S7bijeQ+TjEdCzn9R098Ue/A45S8ZCz1YE7DGdwgxydJ
3KJ/oBEuQX4KRZcP9pUP2JoWpv1vlGkC7sSk2gt8Ee/k6k09WirkGIikBx22bEcmlFr5QtNhnhZV
lVkA6lmob3i03RVTaPPBy0QD/kD5PGSecgaViLFYj7bxrZpkPH8U4fOJ1hqQsxkHBQty8uMwSXuH
TeiQQkmO/gBcZ3KWEQJmhRJTmFfh6tooN0e1dp496DUH01TyXj9QZxYMSFtRpcuIvmiHFs6isabm
GUIPvzrGcuq2FmOrNZTPGKG+FXzRX8JE/fViVscgYIfr8IBozD6vmHYt5zHQk4CbkYeIOVsmJiQO
haHw1VRldU7YpBxVeNio8F/bQKcIvulWzPAj6rnQPh3JV2j4IGEG6wlnrDiyiWyDvA56BBLfxlZA
gLIRK06m08yk7gCQBJTxKCU+6kLn9LYmc/Yp0PRO9oJlnu+7IWqWvH09avtOAGhlbgP0KOyAMMSZ
H+52tXp65fEUxJwQPAv6QA2t6bZOPsIEe6FQTxPyHIpvIZAUoewiiEjJIZ74FA1hiXnW05FHK7tl
ZXffN3pd3UR/O0dZiyAcmzCqWUr6FpuWgHBb9W/E+aVq5OVMgSTqiDrAMtdj4k3XTWvEgvkOCaBl
zqL07Xu5uc9Rim6cLPYiWFvXjYkQDJORJnUIiWH76jvOG1XB/W6uwfENv729NzWdJ4CwIMrPF2cq
anGJepKT85oW7DEWFG7a3xzMPAzxYVuddTfdGQc7Bl6bu7JBJxpvi4ZzdO+j6b/RkawPLLFMLVTo
twQicWWL0Gh0EW/8zo4UT4lm+ZNHoVJpS6qrDpL4DA+LAUZSoxoToXc9s2vRssGUEJfYhieICMl+
Kvl+LcJ9aVr2dLHNCHT+nk88y28iA8XdorO+7MsNeV8obFx3Df6ZUN2JzNVPSOuRJbtRgwMTjFx9
mIkwxEsWV8w+HdZv7V1rFVYpl+i9EQRWuQHzCyCxzWQrw+EtxRrb2uuFa//PTe80u+pDX49nRhZG
4qJDWGvFzHHLEnfAxpmswNvvaH1ffbqtqRl61IGPMidjAbhBka2uCG/IDATDIYaMNTvs/CP935UI
Zrt+pHaf0wYICH0/yAjKJjaMcoFkJ18ToUp5zO89wSGO5ZS6mHt9TJuQQCBI0uFNoUpwNbjVLhj/
UcXOWc692gEK7iaxncdAptFT4+KBy4nL3f7zNbwmUJMQ0kyZOcBM9aFxCl/OCJ6C1+MD4Qb8CH/t
qA3X1B1Y6DeS9Ae+MWRDLdAdZ75PSJjVM7ghGb7olP0EoC+W1A6kzEv4c6X7bbh4gLqBn6McXx0z
D9awM0Zu0TgmYhOoGxap6l1PiYiYSWSbk8N+TCSLPET3o9aVL1mttSxekkcxJbFjYOFapDePKk6+
YJN7w6KsUOYKFGCxFWknAXplzmJtQPp0yoDiUPf5qphZ3vE8r/KqK8u+aaU2S6i11qiEVM/1U/vn
1B7b+vW2hqGdQrB6ufPj02C73/Op6LgALDUH5OdNOD3RokeP6VxheOi3aoQJNgF+nlHISdr0q+9p
aAJp7zOCECmqt7J1/smKphWz0nVS6ypWvEShJEY6S/hi75LrYijSsloC0Deak5dD+lq5X18zPiWS
QJnrirMznPhiJrGs8+non353r0deBGHuI2Jpbsc8h1zjYo5Kc2qlM8LTeFyT9FUyNUeFKeE1oEO2
1oKRa2CUbe2EsXeuAmNLIz7SGcWqBzjeKI/n8m2NRlPDnSU9EDw7Ey4gV6X+qobA8ASUdVVSrZ1V
bgrgZkH4cRze4LaAWRrieeP0o4x/ULKiG2XSRRitPa3wgbVbRkCHzr2aT3jPb6wTxNoDBn4mZTK5
MQZeU+1rrai+uyL/0Um3cvHLVUEyxbRmp5DltKn5ppZgmh6tkg1NkAkTE/4xyICGWV0tojxbrksf
QT/jKI84cziaV1srHG0Cxnp++pE6Y8qLVuSxD4Zta/5bjbVK7CmZ1gD5Ct4aVz9HvYPAO/h/k4tF
Rmu5RWYt08SfotU+ziOgJp07JMfPhY7mKK44EXpDI+hI6rHU2qArcNhf9y+KSHkFFLj4QLcX/B1a
LhnWSoI6/R8TBaUepVYolI2D4grBJLWT0rziPsPT5WbsJGQ/h/ZY5Szv2GYPWevaggKcViIkjMMH
JPCNiGQfrGjeiEHtnXVxL+sSKm0myoPJf4R0taxucROkTwlLeY8ppKAr+WGYku+MaIWjmNZI2ac9
uVr5z9dITp9cw1i2zcvAA4tAN09TUW9cE/BPrRjqQ7tv4B5KRZPyQGskXYNNkH6t4UDOz9m7zsud
dt0yelmRkp2L1DL8mGynsxXydx7eLnnHjTSSJe48XNnsdb1DMf59s/7hZafx/g7eizxnY44aotYV
H/cZ8+l7dYLtjIXCmTwqEPF64IdnFxi+olmHWIloVostIKzScdR/TLpws9Aa6MlbkxtSOomaDl7n
0pSotL/igIB9DO5RqGUF3n0elaQJtvn2Kjisf3R6F6eJ+VHNaO5eLUlzo9LkkhCW9xphLVyiOZ+U
HNFwFHd61ESYXbzQiuHP2ORqGuAW7QYWr9c5wdlzHtnuZ/P6ZrQrEj8PymugRRDdrI24O5wwWrsW
UgvxQI+GtUndB8m+wng3ap9mMfUuGoueEZYm7FgYyWY8tjxXgc3nKtiDs7yZVEF0QRE7WjB2QWHU
X8pP9slue1ayoooV9oejAzzZyuFaN3buEYpcTUJFMIYsVfEQPOSevc0HO11rM5nlQFcIq5ZYG4ok
wy0B6Sx7AY0m36LIUlgUHR8S4qNkQaHzhdGc+T947wJA0wtd7bBXXE/KtHixr5k5KPk01V2v/JNy
SMuGyXQIZJV2KLtcWw9nvs/qhoi4D8WHM5FCjinDmtjh5wtvL/pEQSkfCIUMQYoIxtveTMikan3g
QjnwJXLAgLvVdGPZ8FN9Ajc8hbeYvQXWRivMg9lxYNnKtuQuOwj3cpAKkt5z1LbNBAqvGzGSZGkc
fVqYQxQ6nXH3HEi9ZmXvUrOzpqY9VbmofQJyR6oQpcftM70iyH8tu0LvMyqap7hBgqdcbA8NQ4Jf
kgDOQFmeIUCHnp+cV0WNyKME73U5pH8++b85gcJad9HN6beNGwAkQRNCgGO72fdD9n52KbyY+XhC
ESzXjkViCyMoGnTohOyxS1Timxuak5yZo/DsF/sQCWbAc2sCy2XhRFI/mBVuGTeSo/5QFGlHJfNt
wD72dzyY4WcNgBsqwe6FIyB0VUKBWSh3No6sIQ3LIZo10vsLPoRuMs8a+5kuSTSistLG01kODviU
Dr3ex2jV3r3kRoM9mh80mt9JwGSu7PxL00PLeafDZtLSLdbJ1J9qEDmjp49vf6us5riARwmRCupD
td5lwjrdYFEMnq5d1EDvQiQKH3xZgo1U0aDGrMrcFvE538XTJIEadg1jI8R23AkHj0Lb+f9Rxsfi
5bVorneas2eIdPXF6CG0IQJ4Oe82NtwejFBQJ7ueBCJVMjt1AMg6WjMojPJYLshxMccbELFaMhPg
btzF2wwWmHFM/ymlL5Lwj9qUpJNtlD3MvmNXHr931BD3UM6SSo7RRcSfuAjTzDOMGc9n5ZVC0NzQ
6EPqljGemll8ZcdEuM2J3FW2PhGJzFy8gIkXVyMCyyw9qpkgkUnTw2om+hU3pgFwqbeOqTK5fR3+
VtzR5+b4Ba8DB1q6Ts8BYt2wt8+ZSZRK6HpUQ2+2/bDYIbAjb6fCIOYxXn5LSQIfYcOP1s2pFqMP
m4aH1kiykSv5cIyyPqj8XHfq7coZjv93gzYEJxvYkLYPtpuQzuyEg5/4P9i+ilqw49GQkEEN+ccJ
1kqtkXVHR7sLxzxL87erN3IQh0hHV/Xie+O+QnQGmhNoTbtHxJdfnbRLoc2VRYXCMPq9upXKiJV4
gJ8PYTBYPdzpfQgIU4tdCwrMx0etUO7vnWN9hQOGE3TF51eoOazv3zeIJJiWhk3ySqUV35Nj00mv
3UZ8WbSGq9OUbNZSPmpzAMezT1/2d7kLkBOVMvcj8VkRRMupF1KK7mgK+yaHy4a2CRDDAP+FQnA1
C0KltBc7BfF74CiRQok73mKCXRjcY6oJIVMJY3PDNK2d0lfDT021pBV3eWPT8jOEzAmoUEB4ZV/F
Bh9zGj3/8nM5lctVGd7wwd1w7Oss78gwyPeG/Ig+nsiq5yaOeQxqubxGYNAu0OOb8Sq4U2kMxJUW
Hb8DLLwB5srZy/MgWguFME3GYuRIFkjMGzN2T7QZGOgh1InQA7mGgy/Uy3RJFNdCV1l61XcSSAPD
P5MDtCj/uG2H0B/vzWgDmiF/SlvpqolG44lwPkVth7TYGBysbpPg6Y82Yq7MB9L0/vA6YoMXDkxM
uNN5zA8h3uZGMy50rqgTnaAbTVgTvtB0/CqwVZJFul9OKHWw8vrdi16iXnM67hWG1ivLSj0GTBzd
PR/mebBlN9Ab9LXcZA+/wYPG2AN14rQ32vvuHwNXnjfr03NLDQLQM0zO6Gtg/vD53cf/YIwp2wwL
h9K+O0vvFOG3xQ2/iwhUFSfp3hGZMUJNHyvFVagIAWyJCwtax3MyaqWBek8uak/rsghMbfZLolCf
4FXiqGNDOt8NpXYxzMpIv3rYR5qREyYhq36c6WENh59AuoqDoL3Hlu80lIQRYmsRKqfmo8e/sdGF
ezW2kYHgQN/6Lt/1J71pihmjbasDZpnH52Lq4U1ruARPsnfBikkEtHMQU9GUmwW6zEDo8GY8n+8/
ODbtmE1IqVtu3hK22jt8R7D+6WBHmaWkb+BliVhJGK+iGmuYmSG6APH+QxBFi5pMKrou+Km7hZ+h
injM3biINj3RbxKuK0iPNlCtVPV28IYqpeRVHaUwbHv61wEVMUSwhfqfWfb7tGyCgNO1XhU+YRHF
PmU0WBLYlZxi0WErv92Omj/QpmMZB5v7aP+aCy8pK2csS4Ff+iiwcnBL58I8ir/WwOpHzUs49tmJ
4Hn1AwiTQsNfxgSXpAuq7xhbWAhKd2wtU4hQtRC9GsaD3466tbiVWfHA3YgllBVR8aQAwLNdDOFJ
TFpYl9hynR3OPGcam4oG6DyaPQPHcoqrA+98cDYXUsSanytRVPj9V3dzUKGDHLqj7Q47V9DFbuOM
81rikpyEwFesf9kW/9UlKlyHj3PGZ3+FN7DJULAapgALN+5ows/H0AM7IVZWzER/pg64sKuuYbuV
hVjsl+2RG6mWdDFA9Ejf9zqWpYxJcLza8FyVqsWHFGVRxzvn6Psxa3WaDXCvrbHBprWfDGP2HEwa
L8WqJsEh4zKANSAx1JWwWtcIdsMMw+1VQUXDPiNIMv1dT14qyQzHULx6VS3Ee8EjCx0iPae72ILB
o5g/sY9ryn/yh6VIQAv48xXfpfZpayrGnJwt0VCeQeTJMrIvv0aKmZ94hQcfVaLn/BHLc8aOAW3t
DUl3Bk2vRNO9h8FJOw1ryNSo6lMNGLMjc7VuBuZoFvFsBQfFIzbkbdTHduDVpWLhz5wE8u7ZdS0j
I9t/INtzCVwebZ24cpQZ0tB1LUWoVvEuwTbUfiFMT2zb3Iv3Zhu+a9+qHgKqeXLCSukdnbfb5357
I/ojUoovdDl6uu21RV5xqul1cive4Q8N+vR7WzAypmbGr6KoMM1eRRKs9QxuN5/XlALi9+s0AmKe
NBBGgn30OY3AWqUGJJbdKTswbL31/T+38E+JNNerz0Wr86boWYsjM3Rk3eL0nzUOkZ0YO2LwvREn
wqJJJyfIn4cGiWbp6Nifle7GXrRTPMO7lCJqMpjbgaAXhq/w5mQH49yfaWtFabK8xuxksEPKea2n
SH9Hio1Es4XRZcOqX/VXMOzNsIBHdRhins55zDgNVYCfUIKpvNMImlMCYOd1rLXsQekPNR1+Pcd9
lyUKDojfre0+fBR/y3M8DUmTzpxI6fxXu+RGbY83b8C208zOKSyfexZ7161TPFteXvdEz7blnMb2
W4JkzNYXAniVF4wEBHdie2iQ7mLp+i9anJJcjfPVEO7+5n51NHNNAE608FzBw2FyC4pp96XlyX1N
1UkSnqTzUZL7rRPt4gR6usIgXa9YC/T169kgAy4B8wXk3p6DSQf2b+3MNHLw5RAY1IzPUokeQZKe
7LGCwHpXzsqG34P6kK0iDgNmkrKfNz/+CdLdMmxsjqDyq1ooAZWzZK/wCkZXZihoc6nCXPWwGZhw
1ZYg02kRG+E4RdV7h68B9QFozgW8G3Qb6OvVl8ZJ9+QgGToZXsJ+xnGJCuuHwyaQSK9UiZUa8TDK
29mlmd1DnbrLhxldyl+S/5TwKWl8MbjFBYpUwj5kv868mluV+1ukDJq/KrSOB20JXqxxmNa+A1Dz
6Poe+g/lx2FssE+1tevSKyOUN47L5JbbMHS4lp02o55lNpbOIkWWSOlJAoF/mXgwf+/YrvU425HP
Uw4kGTowlNDh+EJb/iwiMmxtmqZI+wt1NErxj9C9lI8/a/PYpBMIyO7FT+k5tHkXfyFFi+CQ14Fv
7MMB57V2kvftRlw5MFTOcoaXADA/U93B5q2M/kfe8xpdyYOYoPogRnn5aOuoW7bhAg2U4M6zq4dQ
UBcVI1jcjaws80wCLahhHrsf22ZsusAC5eIyPIuFd/IhnWaZYelmVqUWTKkk3espT59vMFXZxqpp
vw/nVISEzYayByXsidnMUI4y9l+ZbpBCI8GvBhnATpu/pfX35SaSzVb5bFCbXwpL89xkIgr5Uf2D
Wkn96jT37x6TkbTAzXyCFzOBmkZUnBHhReEtyIqBb3W6s1sVAlAGtKn38+GIvxO8nVxMWs3eQlFW
48EljEurbJriXacFc+1L94FOBY2Wyc3FYTJneUMHRW+oWAOl+IkUgiAG9DPspSHGT9l/qFKEXZJs
04MuZBViDnoJndYVm1XuZEFluxqlPNV6fwXNoLp7tME+e71764HALorBiAAaq9M9e/XovaDS8i7D
/5PEMHnBKxotmSLWqTi2oHKdBWYcFFLvGJUipvA7+WZrNmEwSwNcKtOyyCEuLZQHSCUO9VJoMAFF
oiTQlQaG+uOJyVGFW5FXj9R99aa6xxaEa4lUfqT9GGB8Gl6endllBMsLFrYNPsT0od+Y+xDr9lg/
AOYodd+TCKZbWxCSQa8EpmYa9BmgVxJyV3gr+0Zy1qekwL9/5402t1XPUzY46xQrsbEImrPsctw2
7ajj619mgbopsHUQ/h+NfFZwaGJKfHNE4LIev/kP75TS5LKGWFojTYi4sJDTAaupyJKv4IWIrMmC
s5+gvAdwf+38R159Is8R6B35RWTItLcRvLxZl4740nocq4KmDBzhSrNy1lP1ejuWB8Eqlt3hxhV0
FU1pCE2iWFJdPEevpu7ml66hDfHghdMY3lLSWYJM+suTAQzpAITPFhPa1yDxnt75RutjF5gNgRXK
0qjDomNPzTawFhYpODL4UHSKsB0uYLU6TEMEzgU5RnFE8PuKu8cfz5s4EB+NdXhNLAAG6UwkQ6pK
TjpQOOrffJ/Oa9/mGdiTxWmFbZrXvKQYKjzyg8oYKQ7TegVkXzSx9XLSP4Y4WuYgx6jFZlFwOQ9f
BB24Jn8WEWxE3jFQT0peKjbP7Xf4EwJ8Wq4hXEKyycOi9WS2VP5TbpajZTTmJ3OKYnvoN/SfDQTp
NUiGJ2mc+xCUpC4WltOPb9K11+x7ygm/8wqZfWav+pcCAEJsy9jYvUbP8QQO5i6QfOxTS4TKJvqG
WhyeaqWxRJdBsg9N4KZg5W/jQoPNdEJ64rq+rbb4i5+VHKB6eVtj4hZ6ON1wGzJsq328OnVNOQC8
vv5CxCxLXm6K/OLgUbk0mdUHZR4kB3DjzGuz69gwIVvd1Hh5BorpDJSsggKJf+elR6G99x4xWwQz
DI4TwjmgT6FEVsOXD/WtQ1Pr0BH9AdoXbB/HogtzyWGpXJSdSKIdfzB5Yr8bXwMAOKgbVewhSv7+
gMSuFG+kXwvkTmec/c1E3TE6RlIkzN35VhXe3dZ2oxmG7upDL5ZHdcWWNz2cFWJSAdisVfSIiRsB
TnycSiMEw05DU0aSChFPxg4OQtv9RttoU9nCrkOAc4s5i/i+fzfa7fmLjbZ1S3DHvVrQiNDO4gqZ
9ff5Qiwcz48l8bzZrdtud3xsPJsq7qG0YhbUY2h7qgbwtNXBpMrUxXXtRBpG5SAJyFe2Ma7siYac
IQveFkhg65aRhwUt6XlyhsQvP0uQcm6n/sejUJK40+/WFgdOfJlvmHEsoj+AKcS7k1kL+U5rmIPM
+j8CMY7YKjbJjboxgHrmcx2eKbToS3fN7tLy8kuxRuu2Edyq1kU9JK+sM8torK7ar0xQeQCk69KA
Nxn/9ofreUTmdS6ohiU9MajXmE6irWhmnjZFA+svn97mq7BkGwWa+6Dc3+GDbpz9/AXUCg9X5JGP
Gshl1Bgz+UzReeqZwDlu77aMdVXR3LKx/0MkINA22/hS41iaWINkiZwtZxvAc52lC9llpVdkyMSL
8g/LdjtU1CrjqFnv24ndk0j0pLsFmuWD2tVTlvVUcjWUvD9QE+yMHyWO28T1ldqTXUUkKwPhCQL4
KK0JR59grClHPmhh6swZhOWRDs3e8pkwWjrU/YQg5VAl6ZfalYbyNU3UheZtUm9T5v2lMBwRMNi8
IwPSgG41E0w+53ev9k7ZTJoo/NjTj4ZO/lSQhUSph+diqFsmbl3Y0l/wyyrsqFrHXL9zBMBVn09S
aBeyBkiKZ6sLZLVF47ZymM3Y0kW+QCvz7DdxP7KWGr+SMjMiyWL6W3Sr8536BwsNbxzzmJ2DKQXg
8eKHOJG9PqSxceUbS1zylPWufWKHWfv/8XaG3RH+pNzMgQ1Bdd2oy3vM2YC+ZljAPhyl2u5tkZhe
e+j1g3TtogBq/eX0JIk0DsdbZ+bHmQsBlJZXbKfwJ3r02FF10UN4wtNAkOxLMDBhcbFMjY5KPJhN
7fC2l4BHdp9/LW2myvlQBCl2SCktndjYTAnUUe5N1mgRmahCLjME17Dk79+94op7WljFzUQVwN8A
xtYF2Sjv5RCauM785w57eVOOvh4filUWuMmv0MoNj/ER4ZVH15jjQLqujVkWBI8unZk4r8MGHZfS
mVliXcZT8XrpzQ0OzPVcw/YmYX2VQw/swA96ZQ7Ee6ZUnev9m8wk2xY/XuammThLPEFaWh3nipg6
eWNhH9gp7Rg1gBQlbTt179hLqsK8D9phNUWLtgoUAIhNKwHmOKVupePySOqQaOaHXP5jeKKpi+WF
c3wRZ27WoFSe+9U2L3d3fjcTIX0BCkigVAoK5GWuBvqkEbKVc4kLFFBlWYyYu0PeuMyGTQ0q4tvd
bZMhuNJkjjcUM7sbC/bLkqzQeAHGg0J74QwVj/dvHa62EnM/mqNWPvkQye9ItqPXmEMhl9cv6GYL
dah/v9iGaxl79BUfPczE0+K3lVhdwWO24aLImRST/7HmBU8XpZV9cYQJHlAwflqjRXuRIaWJFfBY
kR+nIgSjX3XDWXjlFNRfwvX55nCQH8QPR7C4W4YGhw+YELYq9uaQ2vD9DBwc8Mao/V6bqcc1VOUg
W7ISMbYWKms+RMwK21t3w/BFJUc8wdRPzIRnFMrcPIcuObcqNxO89tzocNkv2Q9GeiZOr2NU1e2O
StI0T8HsgBFnROacHvBn3Ak/LwYHs+xHXpm3XVzc7y3Y3/oEtlEsM/wYLnVJUZON1epj0AS0mQih
/ReVrbhhd7JyeoEAzobBbldw3WVweYCUQxsZwBfzuDWkfQcZxZ3YNHdXW6bEjKsm1/3XXcWd6fyZ
fugZ5OYgMFCGvVn65gMvH6gb/LVNkyKMq/ASTVK4BAgYoXqZweY2Emdh/Rqyc5MyhcdR9eDgGk2j
+4AU1p+MfnI1GrjEezfDCB52KJ1lqE7PhZ0RE08l9WfGwpv09/VgaSC7SL8sqDwNEXM28NrKysfh
9M/gkdVQ53jDwrkDio+x2FMelniug35mzG7IE+exwxguZs3zvYihDymDRdY9oCMCg61LKBwlQr3Z
VMnaEFhhYOft9wNHADTRoLNL76bvefnf7w3IMDAfObzdcqR0K3vhxp4pjAyfikMwCb9R/3M8UJ1M
MmLCQ6t+NssUWP3uJNEWQcRA1tvFphtXJDABzLSdLi2qqbH1RiMFn9wx0DB2j7REUg5JTAtXHE2z
9xENaHUzkd/jkjFMOH8vAxkcQC8sgZg2K+Cyxt8bi1qGVRpO6DtpqRP/0BnKlcK1e8kxZiN62o51
jc/neo7QjM7HGvBDZesMhWaK1zlNXOI2ZhHYgJVba4FWrTM0JHaVQ48te5nC3X8l6iXcmrfKQAUo
diLeFsNlfunFGYctOvUaYokhMHLfXsaL4i/Eb1MtpItxkewL1iu/Z9Xt/5rC0AanjpWqf9HUKmZh
1Bm6rzfB69v5YWIb7db7HDsCw+B4czfkHmMN1n/fBVLrczFUnZZmovtP9RkKYgs6tnQCU04w/2ZE
ftmrHfgQFJr9jYLaLH2K9YuUDP7Dnr9SJUMbHt/lzVdnXqf7Ns0O7Sndi6inO7tHLplqFwy10EAu
zXdym1bqbH6sgdIHfoQdWCfi9Zxu1UX7CTfSJ16uzwwuRcLMFbDjPSDUaI60qhxn4cjPI9+elCJW
XKjAyLKxTJ6Eh1lg7LhHWgZ6vIJCqK6A7DwuzEcNR8oZXL9SliQydbbK16TX9iV06RGAlkYowZQU
GRIdVLaXeK7R82xbNQGCF90+eGcJ4Gt/69+ZuhAoujySjlMyIUzMo31Tv37J3t75oDWwnopekvXs
qrCl5beC0K/c839fJLmzIb74LiokvWRr13agShpIaJb0akpGt+I1pldJUL/DVrFrmQjFQ6RZMgCK
rpjc4COeiF6dJDH8Jg6bRrdLYjscWxFqKoD1n/Z+/9Ies4u+GsuQDbw0N/xvkT2zY0GHjkT3VTdX
DaF63Avk2EwDHCerCZqhus4X4Dux92OYbKJTwBFNdmIAPBNG70fYe3mzG639ctnhe4ZQgoa78DMO
zqBl2xuWhXhEhoRC94kMdLy8mqOnDFCGN7UvblM5YF3YgVfdFcyo2lJoj5MyDEgpvWAErVeHUsRX
2v/PqhDkeV0bh/QCSFCx/pTwK7lOrauYOQ5QlOHPUEbQN6QESEZdA18J3iVFfOvJszfUAGlJd+lL
KwSEI4LQskclgh3h3MPYve1Z2YOiv2ag88R2u6ZVH3SAQnU16EOBR/wqeMOKygMWPfydQcbpun8M
XbUf5345zTVKN8PHIvj/iwsl68tIrB+LPAd2BKG+uQ9o7VgPY/opBYt5K7JlmT+CVvOPUyGDbsJM
9GXe0tPxkmklt2WOTffPkial/YomX3jPIW5neOYnptNTXRAGiNSbiPGmnf5IqphJlcU2HGUm8rvn
OejN9PhRVe4UGYYceEqiSG/FTBzNTTozQj+ORlZof2uovRxd2S6kk/D9H10u4vPRCs/YUPTiGt7B
h/gq36FY8MV5WFTKo817OSJmzGD5UgzeTsVjj1PeuYtz6Z/n7NsRu+Z8iYL9Iim4AByrNRvND0GM
vCgASfd5rBsvTgVKUci1wc4vI7YTRXo5fRlXGf6WBy+XG4N4xcxZZalESr2XjYRtShM++PiTUyQ7
v/jg2e1bkWtcr6InwiWUNie+ce+s4kC+iecX+dMcszETbod+YxVw2GjotDpc/bRdE8fl/NzXIsyt
2JTrZ77/SCPC3edKWGEpA4fbTD5r35T6UYeVgJ+2Y672XcMu2RQW5vxKogVmhbc6Nd9oh2joFvUq
lWTDdrRvWd3Cu3Nzc8bH+I8taQ7wIH21vWCCrRD8VkBph2CGpTj+F46YQPGWBaUUSBsOGzucjpyq
WavKMQHznJLnAXq5BagqtSpsm5QzbVrbNx0FZKbr5qhtxd9ExD6kVwETEhIUb8xdEwQ+YUIBbwRA
gMmDg4DTGsEwO9mCntLHMAfzufdJ/AeDIJ56xogrliDwA5bNy2xPpGBjLqzmIcAv6YskOpR6eXgd
tooWVQQjp3PW7Ui2LNFtWy/yWuqycNzQomPMHxhY7wYNM0wspKvWmNGuSYLU7xWymp49v2VM75PR
4PedmOdHK9KJ3e78uNJ8ochTSdmwtdu88JG/3SUGcQo74PL5qB5bbPLO+bYy5mn9IeaRNx1BiFTR
GYD2q42XrAeSVOBOUtPorUBlWScMqpKWH9asJEEvAIX9xZI6wY5tBwBZLRc9WnW0GTTTsf4oesV2
fNre1Cxc3p1ODnIbBhdXL3bTbezQ4yCQ1rq9AllYC98MVl+TBLGWohK4Cl9SWGEuzklQO/94hpCQ
mwC5xnrduDapcbk5WNj+29SupVNv7GwXm+VkWYzj806V3IHAOjChqvjDnEVrRADto0eFpzkny2yj
Wuo5SwqoZn16lGnzaBuyySKVV9fvC+MwQxH7G3CDdJezllmTK3XvDnd4WP3hFlyK8soWO2eSgbBg
18BExtbw4OMzk+Ix/85mMlA0I1Ln+03FG44I3v++RUDM6jGiIIsGIzvurYoMzWhglfGWZGf4e7r1
S4oVqVtkVgzBXqVWu3NOPhhFJouqUUvBAscjs7yBDjA+nlqIB/1/bmRnbh/YgF7rZoad2Nc9G387
Me0cKIqig4VREk8Q19XirnwrFRO7jMGVRQ3OTYBYdOMWBMbWyEHCRnlE/4hJ8/IBnllUrr35IzZo
R6WrpmpALaZgrlwXVLTE22uxTMXopY0Fyp9H1YhopIwJn6kbuBe0HLH+ugeNmjd2nBHhfcfhHUTf
mgpk6rdxGXrOYs9B2kr4P/6QNI42TygctE/wVMn+pKon8q2hnc4f1e5ANQP3SfJpAgJBthnrdd0X
I0Ts7MQyZQ0Da4QovyjbSNElFfO+vDdLshKUREluaNd3rgsWNJlqroy+gz7mGiEYAC3BZaW4Lq6l
BF8eVlLFgqa8FWHM7qX8+Zh3t6vqsz4xVuYveMI4OQ8kskCI3ZtsXhU7vQSnNFtDwCqUkGzZKBFA
+nEcwmjAqA/EKSMGOJHkHe6g95FtbdRJKkhpaifLj14749UpcG/QbSzhCWxRSUrb29QSt92B55az
07ObpSbnvakVYU3221ALVvaPdVPz62XfFf1AaQheRfUr89McS0f+xko/xM7V14AZ3C6BumKsdL1/
acIXPbpxk4pspoOHKkjpBAjuL0z0ZuNV/857CaGLvZ2CIuiQkbRTnIdcZ7k86zfXwMpx5XsDWmDL
XSq0gNXTay1eXVDDK3X1gK85OSiC/mQ1gyHpWO3SLEbwea+VGxilW9agClBK683+V/7cswcqFNYL
g2NhaQw/6gbykfritUUwY9gBs1Lauold4j6S794GVKaSBXpKapZ+hh+HLRV6PU0FNvK1sUjNeur1
TaZUSsbSHU7rUJ6fzsHAZIYgjhW+fUNCcIcoB4bGVC/BI+qzXlByWo/VpP26A62Ms+X0l9nO8hlm
oyPey4epytY2U8XxTA0dOtfE+kXTka2iOqkXb13xP6fKqvCWcFkYexm6KtzDMuf3ADnJxFOKtZIy
/ua3hWx2tl5rKyZlPRDpp4urfRG+p2olKBsgdQULSnNXzioCv6tkWrNnXNpVcDeztzhfEgNDZw7+
dI60wOEp808BGXVdcZJwyFDjMB5xAPKOAgbVc23yMGEkZPbHo13X+RSzIF23PkCYjpHCUMKlGLmU
lgq/OWmxS0dApDQ7cUzGBESlRKcLR3Hk1ZhR3MbxUGQxS4NSbpGf8E1Ck6X5FD9Plnk8CaDIu3nz
7pNshY/pPvgba0ZT0d83GPWYweNYXD+JWlz+e3hCbLYYBe91TIsEIPIdrwZfvvVTn8oOA4Bi5eKE
nrtk08IRjwx8YG+SswrVQW2fuIvMB7bCWQgARwRc1yeqxsqkU5b9I8g4KrYDJNLeR5HJo+qbbNAx
zwTYuGfo6punZghRomAKHSZ8IaAVb1a3fWnvuy70ZOBJ7pKZXqWrXhbV3nwnJ4BANTGy/2ZRZoAH
GP201eHfvWwR1lQwIVUXVg7TyXDrhr4fdWB9rk+PqZRVNkqqC8Wq22QMaRPJtJ+YppU7Yka1Uzbr
Ua0xploQBShGdvSu9h9KNwWndFXshWXRw0UsNfwKlOnwvDaMWkt/XJgQg0ddbpZdyDRhXmiscIzs
rKA33F5IH0xYzS/sfNn+T7YYCBBXrTTqyR5tpVKVnkrOyLbk+COJ9G7xv49YQf77ZiMlM9kx2ZhJ
ca/BzIShcdeYyEqqpplC8kJqg/9E+sPxI/4faXrc1353OuSk0aEqL8Mb+zNFQpLiaTQk6clpowVq
83EihSKUWkhReNr61/hNlXKcAvK8S2nKhUc+w6eJriyp7RD122PLiDDdvTdaUMxD3/zNj5IKdhzK
77njL681L56dDbCltrkmswA+gfDrGdbL6Tsw/DEsqZiiyUnNkjiJ6pc+X+tLVAJQ31qlCn2OKjnF
cAkgQG8cFD3Nh0LRutRm2uAsSIq/L/7KZYBCLzfRVOZGUPWJSD+2Gk34xXg4e+1MUsEq1y+g71pc
68OX7S4xFHSzGveH62VIRmm2rf2H3ozYVmFQETq1GmzbABf5udMsVqEArsO+iJzIWc8zRwNhxQ9u
+E08tXfspegDyr8dq5QQeKYtxM0YrHly8Sm4r/cPeOfCNoKMv1+MVYwJOqsU/+uY4Sqwo6l86YcM
IzGZ25Neudl117wsHnHyo/uzsCcDD0i2BwX7foMdVZcpwO4tQXIIueNvgtx9Z3CEmmVs6K4Y9+tN
/3zvR/xZvyUl64SmPLpxisapuV9Rz/vArpSjUlx+CZ/YjCZdwjgLrujXknoCIrkFBwU1mUfrT7/O
w8dC2aGyoKDAWkM3f1UxYLtUfwcOEtHVvyPeEAMiwd4cFGMDP24VZddMsvZC71pBL9DP59mlVd66
DXdofDPADwdrIbISrv2kU4KBnZblv0kZMzmv4ZmZzeT60rRx/PdS6jKgJ+IlfJoTPCQ+oyPOg1iC
MV0HWl66sv2x8vq22I56jL0JeOxaZC6vJN7rwz80lxoAIUebcAUkuJb4rL8UgK87uGOY7owikWBT
J4rHE6gZ4gq5SJ2LEVE6inU6sU7rrZD5bs5wtZinkJWrM+njlPvJM7eqgnx+KFH3inU2sNOYttcM
/yOrm7JoqGNSEHZ9+/F5i3F6gYvIHCRLerwiLLs4mxkYiz6eMAJbRpkLnNHND3B0XrbmSSdTnAlr
ULu0sNYrPQ7qiYwsivSlU/p5wRvcJusW2ASPY0egkBDJFuEDCWHZC168nDWmcdxn2SCIPtcOCTit
RCx3/FclaR9zsBODgYoa5zexNcgkm7ywYWbJBDPsMKsNdN/Cyg9J7D8j7PwhW984L3beAlYnpZGt
XB9I1MGvVGyleY9wMOpa9O029OH+XEg20VQvNHP7nyH63N05kAdRbfSB/XcOZBlJSvJYGVflJFp0
zufPKQRZgXH++ItTQNOW0vTh4dX7anaMP2tFxKcFgCd5Fgt+mrnwwQTNUivmFdClOPu9RNM4KwLA
aIX2hXpjMsCN/AHdc6jiM7UOHWapxECpTVog56orLCveHv2HsyItrivbuSpo+lafnPkxPWRcFIbd
X3Lo94my0cJRykJ4bnRgoV0pN8QC/AQZNq9G0KOzW2skZT0vL9uT6kWAWD2tN24YJ16S0teTssUN
TdrCH2IWs789TN9ug8lSWKMROeN9diUNSM3LjyeIDgsxORI/YUZSomBjvMA+jgWAWcek9h1cl5N6
VYIZ3NuzjMv6gOCpjohnswFpiaj/hqiR3lmrmwNFjc5udW/wwjPqckRqbpkHBWk/8Ep7hQdIYXBA
GtxH+41yKYyXtLOGbpaIGjnzYNOw2iOoYiVZCnNx/KAVq5cxg4bqQI0Bl0HTPQrrhLDYls3XoC9m
wBpqz+0BiREM2hh66WPbbxur9g+BBt0GdtszrraM9bNv9wgUuz3QEQx1w980lAHkjyLG381DhClN
FKzO2aaq/2p1lLd4PCLr81El/5XqZFNFAsTAe/eHVZE/4GUa/NA9weSyChr+0bCe0OlVqa31Q0jK
5W93JDKyINot6VgzQa3mMGgCp2kJ+/9QrXLBPFwVPrQRs2o+SR7wbkpeWXsBIjkmxdJWVDpNP1En
uqpulnSSsjjJWVOcpWOvuihIuJ3fwbVPR3qfMMcLOeI3yv5jcN4Fbw6FwrcqRWHJ82rsdMIjMPah
LAvR8YFIE0ffQyX+2QrDmOx8JHuiwskJk//vYMmD0llYe8FFgBq5x6tJen6y9ElEMadThLWEM3ap
KHt0jDO3xbUT70s2MZ1JUSHbQCY1VjPok60rQESfB1WTtvsmYTrpUeyyNCvrd+HJj8wBoVqw8QAT
yuvFtSElayrJt+SOgeBo5NwVxeqN9bP6vClM2bNiHuF+eJBgcGPzSCQGMX5PepxCxxRZeX1fxiAD
pjrKGEMCC/7/tpKrudWOYfyNYQFNE01qRmFNDeKoF1ZuhlcYypd64XUhbJ52Al9eIGzUKCnckwxD
tHAflim8yXQRFx7+x9Q1/7WOoaA4KvgfXun8OGY/mg77zSjX8jft4ONUFJKQhqOxemZc/23bOFRS
SPnbvaITORg72AO5kTGGnwNDwEcvwVHBcGEjnmLw9macTiNflln51S53H/UlNng14iA/E5SiXMCe
DattOaWjLyRU/0RviBFvhs2Cct20tO72YtEgor2cm+sn8CCSWaTqvsp2PBW0UllM9hTMwOw8FC6b
etmuNqIm0wtGQ6oJhs3B9aGDnbgQTT8U8kL8DCch//oKrvpU3Rvs7Ptsd4LFCSGsbfG36AJP8OT0
NLr+jm6hLItju05/1PTorL3iNTCV97fw9JsDtsdu+bM2KTU9N1d9iei19wwGSS7ml8Qj/JK8ymfk
dZEmfBoPlGpCsJZHhTgL/3xcTLZrMHKvimhbG7n6nCV6Wyc5e+6sxRgH1yMAAix/vYmtToXZVnXT
CL9M0vENMmEOQ07EeGdA1hLTYVqTWrdL6kdjfoNCT1PpTbSG4IkOklBJN1peAXuxedqZ+PFB6KNK
OSzMW6HEjhLijzA1gdaS05ElTS7Hp/7XdVOgbZhX4ASgd7Iu2qmz30p8HuD9hcH+Tsva6Hpt7tJM
7d47Wy/M25M+AVxhaHqyfX1B68DR9BMyMzNXZYJ+E6H5eooqFF9lWfLSYzuMtH7T6cDT5PbG/Y4t
dOjy5zoClxlLmP79etUUAsBFa8bC/BTkXsip+Ap7YaTHipkHfT3PimaWVN2IRQbdIyT7Z0koZZnY
/C1oaBkHXRMcnyAq46O7icmkYke0PQx6ihQ12pVLgAVVMwO5/6i3VgGNnZbc+M0jNMV8rTusOrbM
igqFlHgZljE4tAGoC+eP9r/FMwlYbSJjIKScqs55hIseyC+zUHtnIDJy+28+UizNsn56HIJypJvQ
PFvW3fP9Givv4MJ97qQfUKd/iwyhz6QJPY2G8IfjCJbDk1OnsYxkxveq6+47tAVUtwkDFXzE5c4n
/G77Zww2tQBmVovNdSBMzTK/6SSvRQFDT6tvNSecTw9oRrvsxx5CNKdb8Qz859aHa4ZhiRnRRCWe
3swBnYxZygTjvrImPmGxKU90WUKrvsCUk7ctkZcV5IN7PfVrVm6+zzL48KAMZd4g34APcWiDMhHK
QCwOl9+YzhMVS236DB2ubSH+39HOLfxgKt0LQlzfLFbJXpCavm6PKUDZZrRT4m0++GTWOC+BcAAn
MtNX25brYqZkoRZ+/PIVsrVQtG3t56T10/rjeHFdAIaXUVEMok02etma0UMPW4CRRbBti/2Rs8GO
lSJxWqqwglGeWIYDrI7BMT9ayFDRHeiSfdQ47c6X1N4Ii7t8GplNHmrb2nXcd851sAZ4qG3SCSYg
wXKpmj3DMlVJJnvBxL/Wmh0Goo2IYvYNRpom8sp3ati9qJgZDdoatjqUB9YqoFkFmtBWI19/v5bw
jhlD0OzUrkdDetKSlD/7wCczH8w1ikZzZSMV4xjBc6GO8EnrK5zI7NYx82uTatuu7/z5Uj518b/Y
S431uUWny/hTrXpYnga72oOtLHtUQID+/HgM3e5njB+NtUVoJLBfca7wVQKRt/8NGHmxkR2z5Rqo
B00vmYsdJzuZRIDzeEk8SQpXD2kQBEMHyOQJZgZ4xMu8kmJ1BMxhZFWLRg7ewaMZWL5JEB0gXbhY
5l1ONOGWNy7+ewG1qS1KI/Sy5+t4FSU49NyZwUshXz8HPG2DG8FkUISlbKc9vX4d8mDDhqkiHGn2
Dt1zO3HIUut6Ac6N7pdqqx6s8CMxa91CiNzIJ56C/dlCT2GYi3eiQOxbgpuf/Q3t/gXGg56KVN0V
PV3gXpy+E0CcLDVZccu7F1usx851BMlbwcf9RXbxUjYGngwV6jGUASGUjZNJa9t8dgKRFQa0p9Ul
SNgBzxNBypPR/o2I3oUzDx0BTTZJ/xMrR0/J7Sfw24mLa7kgO5K76NpT1IqAwF+GcK+vZfa5nqYU
pOVj7yYMmMS/EreaOFy0x32tWsEeqriTekv3SPd1RZJYd+ffAvsYvLmEGUg+HIa0N/eZ65djmiAh
P7b0372coLTgU+/05gP4hZLGtoQrzqpYmq+GrqBZlL4wH9LIPb/fOg3eui0ToidCBpOnDY9VdgGV
AuDBlegzuY4g4upsJmsmjieV223EkWoblrqjlaGtDEcqnogY+Mmvc43HyVbjso8YQaKGOyt/5TvY
tVfi+VoAcHtBVqUeagMwFYXEfYP3l10Tl9DhujlJ/uOvKf7M42iU8zhVNs8F0C2zT6wXk1Uealhp
dbMNNe66DthOqSDwuVdLUijHA15Neb6JxUeLjR40wQbA6CiyfPjKGI7FC1d9B8KFe2nh7nZbdpaI
98JM9pOFbZzlHydxXE8mBk1aOySSyKYmPH2J83vKl0ztUqzJoUHCQVfq+JmNdbFtFNWlqdzf1mge
ti0tD6yqZFxP+fKrpZC6vRutbT0vrIIAIzeFvJLCJcyPS6P7EmywcL7Z1OrwcfKQV522NHHyNYyP
GM49xXDv04FN0OVozYDB5b94/btzp16C+CFSyHzf3SybWvZ99Uw2fXwF5MmIcWj90WwRTJtiDBXC
j/ueLwa6vrau6GW2T7K1ioGyF7ZkGQ2tGTdzmLPCjQgiRwPZIKBrf9O6I8jq3PvY05pgbecnS8GD
HUJ2+mB7JsqZHC2TBtpBUWowUtA8EXlNxlEQtgy8vtdCobku6nDgNkhpQ19302oB25t8Apmb/X0K
PLdkJzu/0bZV7lk/d4Afgmkv57BPBhx360/hB1tWo2G4vrpKDTsHATjugYKa/3SvBZT7cX6CSAnS
FV2JQqKPuSVYCtz8A/bBcHBv2q+xk1iDtSogKXWWVjpm2gGeCQ4kB6nRUK2UOwk1KV2Fzmb01hSM
vmm1/zMrSAEPggFHVYax46Z3pSMpcX8V93M/hRQwF6XeSNRJgacqdFP8kKUrp9/BPgMyTwU5uflf
/me8/U8XQ4pg/lWPnR2EXFm64oRhDhqpVPKwzeLZWL1XVjhRNApCidiR1ikhRIG1sYj4rTnJZPUB
8e8nWyMS8TnTLlENPI189EfY1MZmk/dn5eb+FYqbttfZMcuNZqDDFufMQetEMo5Wa7oJ9xZPF6+D
XKlmalpbM0kAfBC1NK36hbYy5o2sdOiKFcfYQC55839VMdYB1XlFQ/8zd2WMX2dGNcsr1c8Clxn7
H9JYvpT0lbZbOhG9hp/zT/phxbudJphxBl3i3Y5zI+NVzz0ECzw55jkyKoJVvhXBXwjCfzROauGn
pRWkddLWRAEmiJ00oTq8ODUerSPIaPCaBFD4I/ZDjaD1nZja2N66JAmtV67w30H3VbNU+Dn1a66n
vCvvdcE/wwExyVUtT0NoOhEbbru62/OJlDm/rTKpevNvJKlxUu9dkr0twapPAk3qGBOAyv5oTGjt
w/ksEUPazan4skTDbtH1VIoeXCLpISuEAQD2VRWIZaSlfAjlKoKyzEKS2Z+1ioWGjEI+QMUphoLa
tLL3ZAPuNZFIHF4nNdgCzihTUm7eJzt02KJC/AHTTkuU7likBenPlYiNfTlMlxq05QJo4pUAELJA
2oBUzZvIJvvck5vLkiqZKDUUmK0W1zLG3GSZ7++OcLP0LJAEFC+Bg+K2ClhV4tzk/1ZmG9fgetqo
/OO+XUO4Y+ZZgKTzoXuqNnXoxir2LTAinD89CgJaz2tZ1g1ka0Xl2EHfjV+7H8V4r420ZfDOMrZo
TieqrtshU0Gs9D7Lhde9RdCrm9HwBSe6TwSTMJzJzi7OYgnPbv9zkfBF0Kw0sSD8eVKKncW5t0v6
zWRQ0DqfwNSZvAynHj9lZr/G9nng22g8yXBxCNQmuorix/Cf+rlocz2SdouZTEYSadYRCMOuIZyB
fuwOMUsFxYmsRHK6zunZ3zZvwdt1MAiSV2TjuyNbBsI/PUncpi1xgEkU3/vvRPyL5GUC11T+JR4m
Wo9HP31JA0BOIgO2ZOqwqE2Fd0UhO+BSbIP+5kTPllCDx/qNJvU+4srVSZOEd74vWtKa8K97QyuQ
TpPw5TRrT4SxwIFi4z3GD66FWKQGtKdYCXB4c68fmI0gtv2XKXJU+oE5Sczdi/ogxo/zsDrcRFt5
r8nzJexh6gMiexcRLkhoz1vOFDz8j4b5CtVSJ5GFBlPs6OiyLHvebnPKa2YRAH/3RRpsHT1wictB
8krFz2pixoBO8dpxliA234iaemRkNFweFXqkNBGxKMScxQazlzdXbYbupqiqm1aVdSjM1uDNL+tm
VdPio+CnEWMwug2BIjFaYSfOVyw6+OKlFlAH49mkT/+SZKudPDCiMPOeoYEXjruHl2FxcTWiyIMf
XOzXR1O2jwNFDalDk4BTPrTg1gSyS63v/AvWgJYHEWCCDg9H69Dt3vq5gw+D83eKoFkxLGg6KiTd
rWHWXJqLY3dF+U6mF1/KifauBYIkY0NwN274Md5F2a7VcUweMYlWYswxQd+BYBsmtBXinvgaUbIX
G2O779InpwqTsXUvLdMH3nnLItTOr8nonmzWbMj7CriUmcnCbh2+opi+43Yf0pXN29g5NghYGEfK
yOBiA06yES0JNu6J5rseRB4Rgsj4pwTnwtPfcO1XyKqs09lLRWVzBkAbGn11/CDVlsBumeoNNzCh
kanVvHFkU9rPeRYUUNgfR+ssPOQC1ow0oDGt0157WADk/vi860gZcBbQAbF4nPrXwZ8EEPKEY7Ax
lZdSpyEaEzuLqAjICbS/BBYmL3V+03qOkyvPm19P6clZYno72bIyqNcmkrZzgHgrviy8ZhOuXY5F
JN14B3nHqWWcB91wMK1kv+Y9kyeRLR97appo4miud1gz0aVvxqLwb3HKzfAzf6pe4RJnIzr7S4Fc
keT39Zv2QnzyUPCpBa4iAE20NRiJjImYd2I+UJwKupMVzhRvT3vmEI8fsNSHgfWXStJWxZBJ+bv+
VITjOhgRE/Z/zU/jZgi1jmFOn21x9Z+ek0oALiD5lmkKhiEw9SvWC0c3G60OnLgS+KOYagPjnSAu
3R4ETHaE7CQ+yKeGdQRIQ9TDCK/k4MN2ojmMDFT4OTwZ9s5TC+FY/ikvNX7kGO2t6+ZfWVOR4m2X
QcezIrskeWjGwb4wVstPWRVMsRZRy6no7VUOhqLz8Q4joUDBq5FV0tFzfxyU4M6Y4+U4zzvAF6P/
0tjLRHokvrlx8gR8YA5s/b/RQhC7TiNS3QVV+2TpvUzgWjjkVWii6dnzfcrfFVRHktiOKYMCZT14
bTpd37iB9K9dalyA4yIfjwp2oGXRXl1tYXSvDht0anOFD4nEP7HV/w+IsTuhV52lc/mlOq6eFWY7
JWw84g12YWRV/JOkSucf+9rCjsXdxVVNoMWodBLTGLUnUKiEnsv4Mg/Q+YYgdNQWvpvwK4cGQypz
ryeRhkOfay5EWmVH0xokUFMPdWD4zKE6xzanLkrb3Z71Px5T/XxhoYWTqcDrLr2IIbNCNiR0BlnS
tT6Hg7FB4aZ5+QRFCkuQLaZvhjIks1BPhPvQfiTuiW0EShyEhannDtG3QvuSxYuxGqyWBkbwcBa2
7VRGGtv9gIvzwl2PS7JdFMT4E6ZQl319WRo9qhvxlMt9M8hkXHt1MZIZPSXSX2jQmZO4EkCzurrX
2x9f6wWXSgAresheTt+duyIG3G4E5KWzmoRdP4lQ895tHmtiotFf7kQ2rAbIlV9u5aSBahFgKVR2
UclGCKwQrXWfS75Mkzbcy/Np+OWhdKduyRTetzkyEZfTxDLLxp1WaDph2hwTzWw4Tqj/W2ubAsJv
uT6bR7VHOlN0fjck7TRIagA1BqtWO8IEj36xGBXnJ4dp9WKCBKLjRyEHGKIyH+8eVfvtgdrxlMqw
g7/1LZBZk760LGzgBwudB0qQm58UoX4khbbelgf0PHtFF7mzG508/PoPLv8kiShoNJZHVWsgF5O8
9WX1HtQwpCxEaVdx3FdPwHlBIVQv6ZLhNssrT4RjksbcGV+2edsIBAWn25K8YTp9MidGI3wKSCGW
kh68zQcZ73CiMV1CTRZzbeCJNXA98pD5cNr/8bvz7GGF9+VFlY0tlE5ziZ4mOKM/Cel2FZiyvhRc
aaTSq/tPJuLBFOrquIxzgKBMt2w+pUKqS91Jb3ck4Hb6Vc1BUFTY2jBfddR5d4BCN8BqHcgLJnTh
GbWykGdsJ8xT6LnF2qBR0CFKZ6JkU/Y4qfL+uIU6GVdyFgV3Di9gCcpcwLpnF2hQAipDqLAgu65W
WAEloOnUnULS8oMvrNFAh7RMm8WjTas1/yHRVUC1YQfsTk8kPTS6DP5DAtFYKmRikqe4hnxlYAIa
eANozjgJMSGVDY7kP1YyPpii64GHBhkl0gteGsD4BDla+/KH7rAi0xHN+N7/PXbvWU1jZSTfdhD/
1n7c4dBOxVMUqxmB26sRg1btDuUewmVRD61K0MLUEtELdB7fqxga0VWSlNUt1QVeNEqidprsaaj7
LZmpXAl8XbEElDHTFgJceUYqT3mDetsv8ijdLN8XI8+0tHoJ9DXbM9aC2UZJ3zxGIbsK9HrptdTg
Bc3kjKDk1aJOYMnDKvU6CvigTTf2QeSyKMdjWLwhyq4yB6+fbRrhRH33f/1NSO8GZwYeeOlV1WMD
yFtUxhWFSc3a02ry+wXA1nCU/+KHckF7OIovXwhTeYyzpQxhcpaepjff2rCpmzlUbCnK5d8ceFdm
u05HqDbKMtyc/8AUgCDXb3nTUng9MRQTzM0NPE54L0Ra9YXNoQsP410SwJKTYMk4Ta3fmkyLheMR
uQopsJMReW74ebPofuR4k2sqyACaV+tSJ+hipU9HQ8Eb9l+2hL+/O0U1ylfYlI7MX30jVo9PylcE
hntv4RGvqYaOEiC7jkQvMtyynpFlFydNFNmtRAKgslBFRwjiE4+XEHigGgw3OBr1MmXTijxf7lx6
wC972rVIWPQn9f+zLUdIyEdNsg32ULEn04cjNUvWsFnwoBCKQIjkord/8BMomQSi9tA3WNgABl1I
2RWMA6rz5ul2vFXdhqJPbJsc3xnY4JlJ+01kuQLNAP35B5pcoefabRnN/aYuS86Ox+xdB8j7ppu/
Rym080ZAW/47sSMCvlg22qUa4AwxyyhaJ6ODN0+3TNFove9mq7uxmyFxNG1UiMk18FP5Zs2+BATQ
vVgOj+ktyZFFeoaJ6/fykZmj3wQ0aMrYIONRP+SVKKBqbtIYFakrT30tWE7409FMoAuQGNze0OE+
3PdKB4ZwJEE+fUYkR8+BXciQF7Lol1J+RUQYnhFCKtFJe9BB6HYwRBvE+EIooKY2w8R+hg80g3Zg
Le/mghT6MEQ1w1vZcfGTozTWDpszkwA/fF7111liABtVea6R36l/rhvwXzd+HofPmjX7wQplEPCz
yRPIrQWV4QB/j8USIDCz+Be7Fs1UWVFzktwRJAklzgtMgVwpi8qsV7N215myW25k1kDwQcQnxMnc
2sDIglQkmP4aRXqydUSVI62qVehXsxQEUqqF2LoDc0yPTfRsPrtO54F7MiErjxQpwrRvAo/U1po2
d//r/Uhndbe1cblm496kV16UP3cW0BRVINKmN9jpLiHnJJRa8+NqaH41y930CSJbICco6pHc8l7F
yKbpSmH4TqMoMPg3AujSd1ZDhAiOrk5p2E+9DhjMmbw6upQVZSVaptryy15bhJjWgCgCD7wWs9yR
EytYmwR4L1R5vwBlW8dXtdFQAoK/ikORgmUouHk5wDjqsg5MajlbMQqle5DluRMi8sulwyOVaXpC
GatyEoWMprTUvVmAEeOBROJii36xD4H23UOturYEvqRiJUE4ur/t2CIE4WjICtMRvV7Ac96D9f6c
Q6N9fbE5pNYgUA1xlYr42GCZ8tmsx8DBFC0V1DYhxrgwIloRE3E06K4Nvb1Ay3/WttkptDHmarOX
0+GnHJ8NKhVFHy6YPo9NiFH1JtVJd1E0SfPh79wg84HfUPqJ5hMLyc8U556lvDuiicsYfiAD1fI6
TVv+Xs41aKyRwFW8P8TLwXz0s/T2NpSiKs/PFil0rMFtF/YpyfyfyLciwzEvHUCiF8PvX+EWnwmj
WLmYbTMcbteuvmR/UiJ6yGVIEiDdwcKntVdql0NDxWgap5WuKzakmI7DCU0SDLJ9FIZj11F7z0Qu
0ujxf3l74CkwrcU+nZa+PD9NfAk0pQNbtpNrDYQEzI5Ut8NJYPRam7aO62QGUVH1xAS0tPEA3w3e
iRZTBhEs8zmPJIp6+ksTr4zthVQCM4d3VR5g3B9Zra/Z1u7VukLmA3yc+DVftm/F+MJ+FoNjGQFj
c6DN/A/Z6nKtjYtpTi8fI8E8ODKl8PY2hInJuby9z911CVkfwLCn64ttZ1oRh/NEWEwdXD7cq8Ls
SpexfZC3LPW6xDR4XLHJ4oiLetBNUlHzYSLOs6nYKOx6p8+DipyRCtI0E0bB8pawhqPVgl4noYKi
C44/sFd5Q421V0eKXz+s7xMUU+wZHAmsj39FwPFxVOEYK/SlH8V9ZNo5Hp9kC5IB74bcCAOJaKhc
x/5yZkUM5mw8jjjMf4d4V+Gp6/07ysmZ7Jn4ObayFdzY2Wb/8i3Fx4HjPNATERLmeWXG2KXl/5jL
ibUcokt5gPc6wPAJBcZGHFqHFXUDaRVWJ2GWGegg6o7/hJo5q4hs+XODMNwUr+MhlD0KJZ8+1w1p
SAvCWTX43rx/+48bL0PKIMlOwBVmbTdRIU8LyOMMG8/rdXIC8qddSeAf8mIZvyT5B+Klr1fY4yFg
ULxOZnlUeNZc5W9Iq7hdRV4wCEsOU6msVnfPQt5wNNuBY5oBbTMhu8WHRfDcGXXsDBcePNbM42h1
nKiFoz4V52cmZEkgl2pe9HmWj/Ec/t38ljM7dCE9h0s+0M5xg7iNxtrZyT5B6a6K5CogAuAagAnm
BDP8o212ZvQ+cHmXYtiGZwXWCi64zY5OzWMEO27E1tC2Bn4YoZlKTH2IHRfsYaC21pSXSDLkK/6O
iT5/LlgEC2yIf/uiJt6ASWQziLyQTbtPi/blTujOgkNp0VrbTU4I8024fzgtTpnDncZfxld2EWcd
84Hukr/243N0IgOsvCfS6pAcJTC0Ypz7IQLy8Oq9gxFque4aHKMVnL8GBe1qfR4jevK6ADLC42OT
9IICDqmgqMH0mhsZkf3ts1jthxYA+pH+Mw3RIrVMZOSP2MlKJ5ppnkDeiJosos1PBJHVU9CfrlNb
svgsXJSXkg58XVT/GDEPUE4edUhjcAfFqinlnOnOQg6lQ3u5VdMXbPc00GfCmrex+09MvAiwxtUb
wj6eAIdQ+x9QVnosqKsPPDKDnpg+lYxgR6EWZgrZ776TLlRR+p9pdc3R665yLRE78tLJiKAfq61m
1Mxmyc5pOcf/PG6Z59ZDMmga4TsZSeZsqSHyRIMpj6A6fsSkZ3dEwB25R00JRN++T+XiKPw31oy+
IT0hl8Hfqdrr46edBq3SZSIsUhVP1q8SD21Zk6x3rUCe0CdmFHiYyAFXCQ1v3o1C/JtdW++irKZE
wiRmZp3XqSxEXSVtVbNdm4yL0KLuy3FPIs/lHoU9u07N8t8a1kTCtqiho/jvhWz82gMiG0cT21BH
LqN3brdYP2Xugs4tflqqMtUPHUn/uKiajGxI3kVeoEdbMxl/E3l6g5aOHE0h4yT+B+kEwDS/ra5Q
aKMKsUFqiaNtM3K8nUPhMf8PjcpjketP8lZ3WiMPqTfoKgWDkWqg7S8yPx4daLpRxojyxoNnI5k1
XshATODf86TsHf9FNYvyHnekDqzt9e829u3FdqjVmcXTFeySFJCqJNJXry1aN9SOON2BPkF97ol8
7m3BG0Jc4LBPm9dKdrfz2izW1GCYPgI5o/C1hTc/jjZPZLXzitkx3AcG+3tos6DAYufMgOPQaiAH
FDRka1KJ4emvPnvts/VSKaLFTNXxzB7J5Gga8gHe+gNwdRHafES5ulok7um4G43lcLJmC+rAriz9
2FCNQbDNraNMU6JtWvn4OgeYuW9Kb2/e9gj7RrI73auII4CPyJy32TEet+bz6og9hx1N7H1Bn/gL
IY9pziD58BvtJPwnNcnT++Vzs18R31ifugO3WZhKcDUEhKEVrUGntzIyEjX6sK5aILoogtp5q8Jz
Ry21s3IixIdLvIewRycMzRCvMPsKLeItvkIog/RXppnYbxQ9gRuVo8B+XG9qCZP79TSG7PZOZmEL
hfnQNmLBkinaJZlJZccMo7ZUKTRQMT9Kcru/7q9A3kfutl6nTT7FqmbazXAV+iRkXzI4ZRPlm+Xz
DIHJuoKneGFnBY8xUrpF6K3e+Gt2yKVQGVVKiyvX1/zCAfUaRUz5HduDaR4RSEJzXwX7Gt8cFSTh
RDh3CNArwjrDbqn4eQ50p/lBXxoB9te6nCVf7cHn2qagqLfXb9tn7In6Y98Lvjmpd0MwsqC5aace
nUJpkQfz3PnwLwYZPt6/huO1fRf5JvaPmBTZSmkeXvbeZTnte/gxVJaPH/S1i9f+bT5bwQ8w3AMd
dC1VQVa7jzLmQuU6v82vDbDqCyBP+8h9IItmG3r27ar0FvtE9lxg4V0gIBhsjQIX2/1C3HJ2XA8A
ms8pbrGTT2BBMdHYZubqzuYwW6Vo0epyBajvevlPE37qXm87UZCsF6vU1mag1An23unsGH4JWe/R
shtiWzAJ7F11FVZ8LZtPU+rxhGTRM7d75Nw1bpZXb6ECWBRwTvwUaUcG2kPK3IkFBaMMyM2h4ZsF
BxBw4nyB9qz52IG5smwlBq9ZZN0S3iL5XcuPdzy93fMUfRPv3Lt1QSvKlqI9ipXdK/JUh8d9tCUE
sP1O51vkCti8RazBEKaFcixW7ZIA+pgXAatwJ1O2KiNaNDFXdGjPBhan1UMNyh2urJ0SQ25YkXvo
DlIDAljx9iSyxxYe62B693ZH5JXUKDCjHbGfvgIoH/swMCpiHNSv6d5z8QshQl3+t37mOKeZB8Yj
r2lmWZD/0khtRVFwEarAeXalaKvpaPoeThDn4tSH/7kBLHxT+3VXLRrdIeJ5W8bxJP+wnq/jLN5d
RXXXviMC8VD9B5UVMEnSuHGMqGcO3ytK5pYsP/tRVKiDjZVZigfX8bm4oRPJb3qYBn3jsydNAS4b
qRF4dBsuy+typOxJEzd6l/sF8IZe+tF8LY/xyKiSMkNjWYqB71bnRLGH5erk+425QFUH1488PsEL
YqSnyfzZ2F3A2j+tofVjBaDy+F54vYKLvdG6p4nQl4WYGwepWAoQNoXRPTB9yu1666aZ7fdQRg6a
RW3Mz57rRaR3md4394b+8vJu0R7otpWeG3+7aIkvIMva3QvYAMVsbKhsyDZO7l9AoJVGQOB+e04b
qbo3/MhgXg3Cub5X2ulNrK3wbwW2FE6d2iqhdiBD2dkhYIoGVh4hBp4Bs0qwrKVk7Q7PObqSFawn
kcBkCE9fa2XkX0kRJ+z3Ag2Rp4gQHQSjXyc/AbxiExiPKeRBHrGjLPcIAKeyQM7Z3jFMi9plDaDQ
cqm2Pvfov7Zxr5W06op8mBndE1lOGqY9gHkCgMi3JnMeaXWUFk6X4UArm7L5VKdwc00rIwcXe4fv
MrazcX1DmC7E7gvqXTSAkYmXDzbT2WJ6qGOGOMKQ6ptHfq2rHOV3dmhbO+1vkJhrQGBDBWHeTTJh
afgS0A5tRnyV+nb7s9VThgpSgAbt6O2rc4Xs+2cON4wP1iPq2nA5bDHATnSZtaFxQWBlR1rljFCH
OX/9L5BoufKleAl/N6RHXUiiHTPywTYa6JJtyKw1Je4IsmHTR5nJlktPTLNsjFzbUojzvRnte/V6
b7BH40mVc4+cI2PVJNZ/r+XPcCBtr4IBqjgQTItPOfWvTF7417XkGwJsf5HsZRmvaHLIVYu4qXX7
C64LOyIPaaFP0Z6LTS1FUINky9FFUuk584uncKpShWJVQxdfVff2S6fM4XPjd92eXx4FP/97Xwze
0yt1VxhSwVaN4ZR5qceSVIaXsc3cDznNBOSttWwpukh7agaxJEbvVcw9Zg2it8xX4qowy5gWvMqH
92wQb4sPufhsvNeso6lXGq0VG12aL+AQnGq4hKaAn2I+y4CGwFl8zPPrOhu9VwsqG9ssvyy4Cpvz
1ElQws+5rCxrpMX0G2xfz5EV6Fn8pvx1OwLusGdTTzz/WoD5b9zJ4iAjEWRSbnbkN/B+jhlcC4gL
loUFKQs/C36ZnKRyGHWT3IE69alC2e5rd2o1m7Cn8VpOQNYY3ZeZuiY6jZ5oAw8fx0HoW046F6JM
ZjPv7hkihIVYAvwb/id3HlohYFKQSZjHluRUOs6EA3C+LJjeTqRL/WWdjd6wMZC++LLkFu826jb4
asbWl5wtOhetk+96gg12wZhgj5ruNOPSo41AKWvIyNxuZc1PEHh3HbE0I14LS34J4Mn2EXuGEkKW
JJdnvfqEi6ufsYYKYUcnJVd0SwBLCuRTrAAXJ3FFb9Z+vH0K6WpPG6Znl7+iB8ny86nJ0YXksAll
cqp4gMVUrE4UcCR1M8bYbjqebI4PPV6KDxIeAxOarFIiDqxYEqBEmsDYKIKjotr9wx3H53ZTBEOo
D2KpvMo2fMVrtTbocXHpdgjfTaqE6hR1yvBaNTCdOxp2Ddg/oXv/Vs5ne+pYBe3VOsP0skTIxEk2
rVLhffeuVoMjhJjhD7J3pMFjB1O/SK7XN90SAlerdliu/7f3Dpo94CVUmw2AhPnP8DxZVtBeSavU
6PLzNizZSFCKeyaBRba2G/gSJ0tbuGMVyQ1Rzt/aq1E1NAyRFsJ6c8Y2Wjg3TuoGS2D8h3Ex1n93
svgDQLi6SxfVeqjNfU1a0wIQu0FChmj3KvHAO6s6ujXw3hU4isyeZdFpx4OZXfjPGbzv78Dk+8Sm
NlDC4rEXAcAzyfFvV90HFIAlX5Y6xHhAjF/Wq+FhkF3N2fPp5DN7k4NjU0KAYvQyEbPVANJBPWS5
6O7CfwTlakFjg3YvxhNtyqMZEnZoujYReV+8XqKB68zP0ZnUr4SyJgieBDEv9cyCOfMykXovDtwS
w3+Hq+se1S3zVZE44M/E03D/KeI27sxERf8fZakQQuDur8BTlNNfzIuLsiVzQzMtTziA7WJE7NS8
To25jcuPAz3EhyG0oYZh9N1W3m/5gM7mHEyM0mlSYg3117Ymj3hVqiLv6prGCERVs7M1Tpti7Cgt
9fj8eCYLK8SslHnKVP5bvGLrPA6aHGYkOyltVulH0gQlTf4ejSZVaBw8PbQgbO1uDL79/XXH+sXR
C7E5abL7t7hq8yFm5Rp19PPr7in2HbTf5qUaPnMfPJH+fHlFNEc9oILbLP9a+s4ECj3uuQMrEzYz
vMuZvWiMy+RPVQpzvvhR3Lizg5rbXWVObbymSIPmjzFgrGX/ScayzpEMGrMWDGp6f2Z40NRYkIUM
Ht5mvX43fU725Ps8eqoTgqU6yLqnJZFLDC5n6wQOoq51YFseJ7PfyZJ9dWuywk789EPTRxVPFu61
G4MgFk+e3uuhL+9007FhE7QgmWbmb5mGX7pAJKtU4lPKxFbqmxp5yiLrYk9QX2B91gJtaPRHMvkz
k9DAjeh1Tsm1fvF8zysbKtXD7E/adL/ctAJvfwA07EFuh6/I91qXaI4R/1RvPTQlNf06CZ7RIRE8
+UiRat4u2hof8/X5HGTWw66PdCmMwPryk1TR5B2MMoXgHklIsZreL3oWlimWfzIgrb5obewEg6gy
fYHpXi9eba7LoAi8WnZ/xBjswewTheBla9uWiK+uH5QtpxIj6uhyCMLBG6zRCW5lrSxppdN0n/Uy
utOWtMVjUgsq+nmULfu6KlV9OrmS8x7z5MCDtdx4/w+tPR4UsGitYPJSHE9wxoFL0lcd/loFwwTM
jaN2ebh/yNYdW9cuUPzBzwiaZ++YkA2UMTgEmviNKqrZSJNXx+k8l7UZbOdyLSO6hQ28gM+htA6/
UlqdZZ8cB8qgygX0sja8xwH5gwG3t8h0BoC9Y1MYem7KmpCJhX0lzgiDeKB2Z2FxPxr8rTdLV/EV
xf6icJYv+U/HWBheX0wTLV30IRNy2r+QPKBsvd/TS2gbpkr8Azp3PaeZ9XMU7VP2vDgjREFJmWOg
eQUY9h16AhHok40xiEOOYQT60qmlVc9oQagywY6Uqe2P0obsdvMmoEU6XHeE9CCFqAqvx7NK7Vl1
BpQnf+0qmW4V9ElaU8MSFmj5ZhducWAypTycNrV/WDg/FCq/MsQMTd2IBU40eJvDNXUi9DKDdLN7
Zfa3wruuC3DkCjiAlnNEHemFd265rT3oyyQDbJAFhjCJL9gwI+NQGixgys7jh+o2pGunDV6YfUqd
AT5kvbF256GSHtgmpIEa4Axsb0sEl9Zdar78LDEpNd/rMFEQprDVCuncamlRi4FWYALtC4bsCbsw
BO1YG8RH780mZ2sW8EdkHlB8P1ZDaFTVg1UX7oHDh1u2SIrXzyKaQN2rW9uAKzxK2dnpbtLpoS0a
5xs0e3X8zc+YA/pYU8Rnown8jR6c3ZRd4R1EbAx+2uff4ruB4yhViq8PyTs9W+evIvp6Qz0WMdiK
YWJwT83qHvUeP2KOzt9xWXnFGy0UDNG1UBFxC0tCKar+CLlkVPxUIqs55kFAtF3s1kC72vwb7KSH
K5GMJqiBrzkXbmBA3w4u+kUdbvzp6A67W4VnpxEai1MkqAhFPPsCR6Tl5t0PifxSMAxBd0kbX+Qz
hnNqvXLti3mztMV9wMb2jiV4HAzFZbuQCjD6Y++tfR7IuShV1QAuOhpPyH3DNcOX05DR+eZLATXD
Jk/MJtxB+qdYW367JKo+PvkGtUeoHLUwgAuaj4bIfulD6uklYqzu9YIpBY09ZRBthSpAXiOazdat
PNxyb0hH+hKWSpcuM+om8QXgCWZlS+ZtXPpQvmENN5qYz4NjaIiO0zAPDW1XCT8CAzYWjh9r4ru6
xc/nOnL30ldnWN0/s6OH4kpFTB0yXHlhpGmSYfve+6luKQc2qvwgF+9wHw3V4Ebb/Ou7oh3sBH60
CFM9ybRrCbenCqTN988T/0FqCScPuCRP/NpFGXjl+1F0GfywNMZo72wQoRjMT0SqHxDjicWLnpTI
gkPvfnsTpo3xxEgrn1dQrBrV/SsxIr3EXNKFVKUzxS11gkVPusX1i5c60WY+yjssGHAdx1e4qFk2
yBagY+j9qhZJ/IdyQ/Vx23Yn9wXBbcNWxn8cLoYY6FLeh7D7mog2IA6q9eUMAce1H4kWrGm3so2n
vnoYfG6aajJ6sI4NuBRTiSH9h74cprZtes082Qnud3ej4bbWNQKTw3b56gujjoCtl0jsHgSkYB9C
ljqLMXxe7HelB/uz4ROkPYm6gqOHWwq6Jkza553KWy70JFwFOWW85I5x9O9VXS04xtXWZOTPYvK3
fG0JYLyOeVd/UdcyjHP+ShszFr3DYgB/IjJqJWE5DoZGroGhLwVHwuci+RCqY98f9qA9Ei/+v8bA
F7wQjwOV3VxviMC4Ib1AHyIfMwMoimbSshxnkeEoy+CdhoRjj2d1qdppYPZguy65awstEXm+xql6
J/rNkCTg4MFQWVxPTNOWhIq9HmVlc7SorDVJsGXvd0mNIBqcSTbzek0w034A5Z+WAPD3NtSrAdUk
si0WDr4UAhgsvDHX8XbdSmJmtCGATYSKCK31vLyq3odJ+mUSr7xbp1RpBDjJJNjzcIr9Ce/dtm5z
+Q7+iRQvNZXFTmJb3ukVaeJvaS94IsrXhAtAw/NYie507k++d0O3IEJyJzp45CUMWQz3mKbVen9z
jlD4GHJPG7ndgs/g3jEJP+PbdVj4NlfgFDmHI6jZuEQYPLDKacbpXUR0WSwcye7WoOMvbhnRI5zD
4nrQxGL5X+D/mivTO9RQEEn+J5+mwo9Gqtba6VIMqXtFkRxpPbsukGktJS3HMbD4qvB0tn5ZsZf9
UjS/3l5unU94jzGWRr5Bxevn70MW70VOA4XL7kdCCGeVE0KhCxVZVIy+zZLGy6fezIJmLL2a6CtM
JM41U/tTJsLjHP7OEsTz5Q/l1GRpI7y6ohWq9jGP4cEtN2Z4SJkCPWrQRVlKrFbW6nSk8BQKgTf1
BGDyTSNv7JhogA7pxGTmgD4OPm9TgKcFWTFPV6THWjsfNGYt+ieAx86RbwY0pJFeETJ/eEcfVL1L
xY6zveCb7tXCvpEdVjGgSS6oQ6R20SDH/5M3yitsbkey1aGRdx/DWt2j+hBfDDwHaWik5LMhyVjZ
Ac96vQSVpVksqyZXzE/qKQlb3LsecccTCDUz+N+wRaNPHyeQycZL7PxKV9r1IjLgc87MKwbpg7UB
l2NMsbT1pzZ/Lk5mC8VaqCy4mJWagZQGQHX18FIHFYTnG40KAmtdssyrsLptQBgnhvhsPbi+8lHT
QOIys0lMBK6X8cShrdahubg9d0jYloIln/XEJE/VVN9X3R5G9adDxuoYEcJxJL1RaYZjVBoUlWS1
u2wg3LjhpSeXQmjMFOfbEp+mAWOL+nI2JmVgZ7FOegMVVzH5QBEeP4OKlHHdN+GDXnsRWRHtcXJZ
+kqgVMspE5MTtbW2kjT5db2U16tK2mvAN0B4PGqMbAziQfJhPMEk+eLR3lN6TCG1aBKZYN/3NO/s
6re9RZh5HwhTTvMJxdVcB6WZdaSE1eMMf7R2BR9A2ATloYwa+ZXMOTxMXcCA5FbKUuU4XUgzM/ip
RhpkHrDKdjuja2OEwaujQ9XNZDMz0ihgqOxK8qPPpelTMRudxKQrT7h0sTPpI63HALYA5Xx1MoyN
k+c+/1+S8xdYRuxJY1R9nSY7Wk9nSSdla0m5P81vsBWM9TRt/s5g0lftQhldFXUg6EVuSdnAWxPq
O/cuEL6Ozi7E4mlx0pYu/rl2NnPVjylSVn9kRPiRTCXLI0hGtqHHgcA72OyziMtq26bJ9YqoYJOM
FJg6eH6eQuNQdAcF2saOW/P3yXmsljK8sbsgoAMBmLHrBsLjDEQQBT9mp6Vjrk7iBFO8AG8grHpJ
p+3hstmY+GvgBM6zGBen9mta8yUB72jq/2j30tEUrJ0Ls3iMhEgh3QS5ueNajzcSWyVT84HspiKs
C/CPCAx9W3gKYybux2UsNLKvIsNx+FmHhnkG4S25/D7ggAYnL12sG4GqnWo3WHqGwEZ/gLou04D3
HMgF5SQWuev5M+we6nNZ3xGsi6Y+JsheEoOxhbu4fDxldp0WgS69r78z4uTOmHEuCHA8Whewo9Nc
SGH82jVy4mWpDfp9G6Z9J6dmwWyCgFhEdI4JVpAEjtwFTCopUkyFIFgFuGnbXH6exHuow6iUHRYN
gcF7RYJkM68sx3MWMuGOKKBNWy5tR3KWf9vXcDngFBtnsRVf7vZa8cVLNf7LyNu+UUU0JJpFdoAT
PWefzkqPIVQV8d2N/7Ss48i+9J5B5erq7tLnDGFU1mgACF7ORc3O+RwG2wJA78x73RxqHTueoCPB
FIWipOT53FgZ+vYzYfqd2mivIHJjkOKGenWfWuBx8DdAp3QWeuZpIseIFfR00pw0ZAQCdJv8hLw7
w8D185HfQCq7PmH3X5FReT8A0zYbxYXxmn6AVAa4IGuhHHr4fJjDJp26+hFrw3TCbKe0p610gyJW
aIfBJyRlcoJ1NmMoUiEH7an85DXM7pUEdIhwJrsQmp9l5t/Lw1MSii7vl3juX2pOQxXY8kh+ryHO
tmK2VbEn6CTRIJlP1tAXnLI5gb7HJXv6HZjEc4K4ArPSNIpiUuSSYACGArtlDsHa7haVkzKZIucL
9o7Vy9MBUDNY4Zg0SX42tr5bvyC85MwuHEeBVE7zuZbnyFmeVPYRsKyDvivgWXh1Cc7CUXoQUdVf
41p8sYq/DgWiQGavtMYSqzYbejSYiP1ypZT/oluXTBEVj5TO22+a7SLuLMBGX81BQbU5nJGFCIcN
MIZIQn2zMhIUkfz1AzEuArEIVG+vQz5frobd68ozcpztcoT9U1yY7F2j93qsCkVnvZELaPhREDTM
B+7HNGv/gP6nhKfvFzsx1jOnB+uFghxPMR4i/RBCv+QQbFMAXDgTpfytP7n1wyHJFvFYxZQB9GsE
+SHS4L4PHXm6qGpygeBqtE4VKT7QK0dRzgcDD9NVrBL1I+y3TX35H1NF2MkBrYx30C+pMSGkytXt
tLpV3tn3xP2lDkK+slPDvGUzL56hdAo+yMSmndtIcACIF7uE9MkF6qh4ktHbsDeN4YTDpXZLc4YR
zB5hNwX3x24JMvm0pEhe4ORVFLSkkmfQTr9uXEhFfpjrKpfYTVL8pmd9vcZcCKE6oMBmJk3Sm0f+
jrhbZlheSJVjGeI0SW6UrcM/k6SJqSAsOs6522WV79F7aK6psYa+mqtq3xHj51G2wPNgdv4Wt5Ku
TZJfqLtYBLiambOgKdsUD/8vrSPeII9DeUO0opnYdyQMzwVG50MibT8ia3DHg/C1oFiYf6FvxWK4
xwkuOCvwduf2Uom40MY447BjJFn71DgpH2CnQgEUSYUN8GNAUWWMw6UTTVZrpWr7qSKrt9OQb5EV
hYHaNi3aQDjz8kLwQO7cyBEn/egQF30LvVAxlFbxeTBKDiZjDasrAN39u/lXJDc62TVBmdTAmuTE
XH+VtGLQcLPNFu/x8HH4zj5oBfZikllwZCp7Ls68EG5hNjzJzfRvs7JFjAMrNIWAY9+Tjxm8IZK0
mNoGMAgNpk7Kb45TMItJeKXng6eqdo3R2bYgOOW3Qn5uoFmvKEgGPSDjjGOd5hPHL6Uh1cs7CW73
rec4RGuYqFAOEMOatBCV/vhHBF6QcPB2prEfix5C7NJhWih/pYvdU9Q37w9kKYHV8xzwwOyPGjxP
w7qGVdhCHomvpizsB0hGP9M48jDnHNlSzR5HzrNUnnh1wRiAwRlo8GWDojH32bQu6oF7KbMQ6sZ4
SwEtJ0CaGs5s6HU0ZHhzvoYM1zAjUwgKBuiql4QVB7pdF2p63Sp/9YMBclrZ0xv8k1Qluvm/zSGo
dXQAI1z1COpwuiHzQPDR/of81u6wxeouF2N8eo4TTcB/M7y5MxrUU8Ft/2/a8xVGaaelylb1JnAh
cZZ1mDZ6JXXDBhkQaGOWmq961JELOPCzIJnEj1eJWsJJ3DgMIuobZ7U5GXSWhXfndBqY4Cpj7J4F
kl6IyGJ8YDkEGsqUH+dPvPQ1T2/ghnRBLCoP0tc0bJGwWjYINFPaeLCHsjk85pEtRM/oSoVfmGTO
1bx8g3cTcxDHQ3RJkSg+nCjuUDZgbpT913TPeTpjJDfw2fMK4pwZwMNtsgkO24JzykeHrOEExnFr
h8kE7bZsjoMbJ5d8Kk6usKDbTCAyU8cYHRGn1/SiNutBfwYGI03UNnbWzkA0wWwBkPxY5T7ZIq+d
wSw4R+ki40EqCigNiSNBNpbm+kmfWFRUqnuvMFiLduKBJF4G6p1RSK5630pln7sAYx9Se/u+GNLf
wLh410jNtsj5cjkAHl5IrInYLK5GdNymBp9Nxz8Phok77rScjTidJzeMLXvt31lVR65i2gudLd3p
mFKmZa5/woBBW+WVRwQJvWseyMzu9b4Dsmkgm2s39k+d+krEb8EfQJ/RV7mOAjPRNiHPt0on5gCH
/Tc77f7GVbx8ofsWXbFiIILR+1FQSTBiXp+s3g+fExPRf/IIFFCGL5pJeg2csATevtWeKqYIMew8
NU/ZA0IX8JhgHicwQEHw/f2AUXE7WTKK8jEU2HWiMUVniD5P1oTENmo1THVnuDTrrTlg1CxGP7qC
7cvPTIIcsPeUA63jHUPZgrKKPt/KaQ0j7XXpFand+PqT+L4qcEMrm44Dovi4Z0M7ZVG5nJzC8WdD
PYtRS7LQErBL/VMqJrEPtwx7fX/sr1PeVQ6MY6Ww2+n+W2dMroFIU1FCjWEiCfGRVuLQYCuWQxpf
vKyWN2IsB7/wgJvsHbRrwNUDWPhfQXH76R4zk9UAHwcbWAheA22RJU+UlijM9XDXNshSPvrIcutA
6f5zDrTRs9V7bu3ZRsR+0vSUVtTfc/mYRl38qX0+dKtKYCZKfjJTpa0izG0kSuHgMy/nlJ2B5YyP
wIHeSWO5rYO9GloQ7BCgnSvwm/98DF6cfgmJvd3A749wfMm+5FZVTWTvtfP1KjjKW/AC+L+q701A
c9PGwwz12WI2+DJQW/mJANDx6sPTwlru0qiX36JFhieJZd4JBEbfsh8ifTxGSvRdhBJ1tJZjllr+
4en1gZUsE2Nau2AxhZVK2tvL4zJl4wd4Mb6x8depcDGHOvo9qLtKgtHqoTAxKaszH10VoW/uERZp
C3y/+xnwoJJbmnWkEBEQw1mG4DhE3/Z4aHzZOOtKC8oWfAcf8YNXePSD9CwZ/X0+jHu7KdFPa6nW
Sg6h6PEVnXHuT4Bk3kCDXOMi6mUnI0lkp8SbBk6IJz0VX0XXG+5LNTNTsxU2Jy9KQ8zoMM5JHjbi
ZSfFC4d1MzJyoEhqz7Js2olNT+V5jGTCBgfbDZbT5X9Pnm1Hund00KovISV9yGDSIVq9xbKJPce7
LcAkPBMTMmUTqUcKkZD8U9MgxbBeg6f/eyp1DkTIryupgWLj/2V9UZow73hhXhKFn2ZoUVl0uGnA
uGVzwxlmWXydG5L57ObQmJy/ZDcDAwPNJvEVfouxI5R0lvbjPYPcqUy3LNLxJoPXdR+A+UmqrZBO
4ab4t6YEagN1h0Ox+ohwZWiYAmG6uAG1ZphnZfQ/bQIYaJKLmwcxCRG6m+kuNZXm2MZ9MfsBFsYG
jXq55Kifhmtefp0j4dtw1q8VOqzR9e5dxY/vVcHN7GhGXYw6KQ3vtUXbUSvJT+Y0nN37lSB9PZzN
e6mmZ0sZebnpLn2D+Ei0y5rBnjGrk3LmjlPipW2VdYeIXY2cTbKnTNbRJOwlZXpUbFFP0IrCudiJ
eNO3y2nOKZVeSqIYyACQi6fqO+Ibloc0UgoFLGfSpWK27AhNXYeEo35DPEKiGQoo3/oO4qqWQwoK
GA23CDOCtMjL3WfMPrjlwHt6Lx/g4JEplua0s1gymfzwnAqMHwxg5p8L6oX2mRzTNbSh4ozMFIDj
g2y3slOT3z94lyzMvi+w5zGM8M8FXhRgkK+X+sGGBg+jeppa5CCGpdG4n21v4thsOMsMa8IQmAml
1qqFtP9mjJ98JM0ZvtNOHsx25//Wr02ffjCVNKZvybNULrFGDyI0XTOiO2uKUp5ZNHNE8kwhe4TP
7WR8yVByRL+k8KtlTUsS8CTTBAII2uC0a2Tk1Q0zZG79u1ac87OZX32/QD3Zkz4DeXptTPuDJ00c
60QiqOHm1+nf1UdOzP/v8z8tvIw+MfizngA8FpyADfjjP8iltbvWR2EZrBN01d/17gMGT9iTzFqk
9vcieJ4o+sJ9/szF1mM8eJ7e3zSCcoTimpgc78lRd5Zxyc7zskZkdxvNxyQtGfJd9SJxWpOlDgkG
CjhSrjxJDOfYIO5cOExlZrhWS2yXeesBR605VGmvL/liF2iKx2BjlBafLFRIt/qJ0fy/F4ADFFvV
ziCtMU44R5ie2JrQuU0qJtkxKeg6CPRMF5G0aRfzBtEfDUP3tmzmeQRoAjLsG5sVqnpxSg2OuY71
CoWmvC6StUqNkt02J++Lv7/HO8vHLCf3drQjJ6giEKBvhyBycAKbCHVNB8HGzHno2YaFo5nGXdmr
v+ys06G7v43HrCQ96xwUxbZ2wulYh8/oAUV07t/57+97vbZ1ooGqhXlXMZypIyIXFuTkx75BOCCt
ccfLb/3co/DkDiT5zZ78KjHa6Bizoje1MRjIAKU8YMmqjmEjkyoDeW1Qus2jH2MoKId9l387dZwj
alpFwi9gT3vLNSBdnGhYpHZuTjn70OX6LbL07bC9RXXuTAl9BcirQ2bWXxjDoNJHTUw2i2bwvEjm
xUuJHdsyuv0GF+qL32/cFFWTRIOJDT0l7JIoE/WZ4B47k3/LloUBi6P2gAR1BKop7k/Ee/bJyo0J
s5GBICPAAbznSI+kIFrDy2T0/mc4elPADluKroE75TE83rSp4D9jBDe4NRmVPHO2Qg0UvsTybNam
7X/S7gE8kvvXHV+5qTKSrsTzDOpYRoxm4Dx2hsZpe6A74l7JHAICh6rxNlj2DxXsSVF0FeYxa34b
uILo/Iz07Y5XMR/XJpfo/nQBW2Egp5DGFylTBM8Y/a7rMEMXfjMljnQdRRic3CWR5/Foxkk1yulh
UcVHtHOKVbGFM/l7olQ9+UKGYca7Te08auDYygZZT59w4FoVvnEKKKHZycDB1I7JsqHX29mFeJkR
W5RPIT/He/ahFsgmYTUjIMrmlgCA3dvr1ddXwqSJGo9sOmRaiziSWbuknGNNzG0eRL+V/2KYDySP
vHi57haIYrwvPlsW0UJrkbgfbxjfLmoOnv0xcPlQnmUukJbxcF2f5x4FPGcDJTMRf0rjvq1iqKj1
8anz1kIpUcLDbyr7qUFCV6MSGdrx+BJm0lvW3/VaTtv/ovpYLvUIweaI3pvFYl/WVpTgY+WKD6AA
g/4ORBBBKHlSkmWX32k6/jhTgDqvY27/6Z+TG0IQRURw5fkLRlDY2CDw+1lVE2gnaoohNwjlNkgJ
T62HaofD6yljVYGpOSO11FcWdK7CzUf5UFbhCmBVkAey2kqdL/pJ3IzAELxeXWjJXznJw7kjrb1f
SJpKegIevJxZiI42ShCKxQh75/FXwJC9ey3fYc4L58Phv7LJWBx8VPC7YA3uJNWSBBhyndgTA6+P
SQadklunpUVMYgn/xB4PXdprQFBjfkCWk4uN+DqurEYye4YLa0dELjAB6HvftW3vQ/lUiprR2DgJ
KKvbajFEzEfidRYVrxOlInPrivO+tAIDFjvsks49Dc7ECas95hBjA8/PB3uXZK9fflosK+8JniMm
vyoYLx2vcdm0zt7KdC+2I5CZMOPeSLQarory1MsBLaXFx5aFS3NEsbnLbBCMTY7f4cBJSJUBM36E
JZNEza1Ef5Eeh+rLUwtqGdeVKU2754+4aXaX074YgAOdqMF3BhCqUmZ8umKv0Oh/WuthUuMlnu68
0y98JXRxOSFcTsVt8gpMybMtG00AlXzQwZYVLYUnRN3Bh4/ZHiodTj5pLRxKsvfKZ92pmvUbINyV
Ti9LSIjhemrH5hUm5zfyWdMWohu/M8YQDaQ16xcH+pRIEvWmHJ6laz6gcRKbpkcmand2kkYfye/v
N+zwgm5U6GGJqwC2rw1f95qTFGAutVVDd3WAXGsw0GuPWsrwpd7fExQwYSB1Bezo7CJchecvPFq6
yiRWWX7L0jnvmtxKW5AbjAAegONLhJSS6r0Tp/3REnt7KuS9uxQpr5KeFlrWb3pjKkb1QnG8ei4y
JxMAJf8SkT//iLputWhfj2VtzKUYzysK/+Zthfad82EiapeaNkhDkVsCdudM5EMLrbmzwGL4dX5I
0N0UoFRKFRW1bn6LdsD7SA3LRRI/TvR+TaP/6maKeX8QBFUUJ6kyn5hkp5v4Vk0VmitEbmOw3a63
u7czrHXUUcvtEy+c6qSdgFUVxxVRTaUKWQTobGSuihlZFYx90+Uu/btK8AOfJFEsk52RIRiVW/BH
l5MqBw2CeSrjOe5wTmjq1mLG6vnBP2w0oconh2rUkGPvOCV6c/Y03PoBUQc39kalbt6ngKnPtZKu
eCcuqWitt6VdbwORXjOo0cnuob3RZwms/LKdcNupi/IVXDQIgwXk/t8wx+SJ1tBZA0FwBSVENF9o
1wjEYjYbaSAe1+Z30XGX4k2kpprTGiQOSTtd82/7zGrQSimHf8L14KqUTJ2l5YhLw6Njs6kc2PJp
CcLSkCb1+bbkEPpP0waI0YcNFozSurEIrKgpssPF49ijZrYB5ZJvDcEpmiqvnhhdNB8KkGptUEY6
bNSfvi9z02wS6ZGCUOs8k4UUiz5Ojhz/ynkTXBGP7kNP+XSP9LV1goZDfli0XUseyWiBCDoaiRYY
PDY7xmw3i7cHo0tivWq5M08A4y2BgFF1ZaK/+adh22VNh4Ky/umY9/5UQq1ydIcCadaUpPzU64Fy
biGa4LhQThxDUtAbSvNWlJVeBlzoOpXvjKDzfIN6AGLziZ0mxDvbIH4We76eMCi/RNKGgmbb8ZpW
cx3xFHQ0/hwpq4CjPW0jZalaJnzRW4ORlKdCc7BiPEcA5cKlh57tbpAuh9pI257qe0dld2Zwsg85
PH4nYG+pcKnXmtQhHejCR9hU4JVJjVdmFrjQvNNM+WOJQUvoZ4sPchEG/jC/JKQWEdfqiHCuaTzP
6dcQiDMK2dq5Mo91BCUjejGAfWoYcN/zcMWlKoTiO8v5VnPw8jhkEd0Ar8SHA0X6lZkCSf93e1uP
mE6+oLtqG4XSpWSB6o/NsGza9DbkyH6H+HMTP2/WZ8nS0GjMV9hDfCHHUMV1QVsysANIjwiLN4PA
hHdDIgzL21MFixAMcYkXZ5cBZwGmzqBdV2FJY68CO6Yt5vrUarzf8Ti2HDNXDy3RbY88oj/xyZpU
0mTK3hmm4YR35D5qVrv0Um2RnjszwCj27wtnZYBgdQfsRzb+p2m6edBlzm+lQCD5wzpshIqyf/Tn
u+cpIs/ZkVGlVeJ2BcQrTiEX0YWt5D+TytrpsRvN9XCu9c9qG3qbveJj4siYXYhQk5U1MjYKXw+4
rBOYFVHRKsR96F9k5PWhoQIG9tUXtnAXh9OMTt8jguNedbwVUaDRix5xYzUOBlbD3Dr4peIG2Y/D
0FzKqC7deMHqcJVtbSF+0WkTXQgEqSATv+egIuvp7+rXd7G3s4XTi7sS9HedGkI13IWMnN/X3rOs
Rr4guUjSpkeut1sv+LoqbijUeCaAwJSC9flWdlsIvyCMaZBoTEpDZ7IcjW0IqawYk8lPL0Y3VHq4
HFb7NdFbQjFqgcP8QttFoGRU++OMXv8UA/OgqsLSRCRWoDe3cg6ZerWkGgmRp7QyLgqn2BTfUUre
+jlSMrGPuYNql+IvcqWxSKbJhWS4okWozL0ITwTXd+26tk/BBgeL/GYxHuLg7usL/2Fi6dweh88C
FNDxi02uQaDgmFhbJG/+mqn6ov14TWMpfAKngfWG+uwPAN4CgX8SMS2lDUF7qRf4zOd23TIuP69p
vSsrJm2XfGgCzeCTgL54KcV+b137IXwDLguIIVwWHVk0zSr6xgcQllb/nfIaHLAKjbl5nl54srk1
Ss36oY8ObGMctmrA8RHWNyo4mmEXrJq3NyTOJW4mLARmdt1NCiPFzn0AUwvgymp+pvCX830ElpRQ
lrw7BM1sC0FM39G8YkIzu3jrpCiE58+A1xJ2ypFQ2nAtApWwb4RawLlbSgceQbcM/OOsB4lO1KfY
5P94o9mh4ExRphgxxJc0A0MsJZdtiUtcSpSpGbMmfAcOy5hbMYmXke4XKKONAkwl5AnhC7mtplkT
MW5DLrjWV8VPSbN/o/91rr0wnK2VOccztcOkN14bHzPvfttlReREGHOBfLsx+RN/ATZ6Jj/hZ75e
ECLgNnPSeRzvXIhV/9OPNfD4seC3qQwouvSooc/oMArA4laqTkv4QkB/IxRE9LRKj2Q9BgJ2qQfG
ju43wZ9Aq752xbdwUx35JUS2B0HDOxOcK3/xk34RhGCn66ll3PPwj7syq42xxliJtSDPqaMSavEX
H9LTTROdD5FI/ElYJZNcC7E7ljZws3Da5vJzv68+3+P/kbcNkm3K2eXzp10/n+xiL1GZ50UA61rc
uEAa/LQz+ae9ybXM4d6ZebqsnZshx2+ecIX2XuX98rCbMj3rVq7NUJbicbP+/5pyxHUXWUOl5x3H
Mep8oScZXrMbNIyk2+Rncx2uVneg6sXlttOeQFgeoxBbkR1ScVmDH/ZX7aYSaUymORI6IGoQbXBI
uFp3rKsv9/Opvx8XXgObKDCrhQN9Z5A25dOv0frivHsORmsHYXduqTOyFY8mvDbCzNcdNvBIUi3L
Tt4FlimjkNTii0DJyhq31H4j0MFuR+GleFgMPq9MlCZvB8R42zJqb+qiv8kpsFopY61oBj7mgkjS
NFIIGTvtxJ8c8L8bn3n3Cwfwqu/IDX6eGKHsKmae0+U52LR74cDAobVs8sgdP5jdJa7xWi0BfNQJ
A5gZfJnAjcZCapjI/kKDXEVe9PrTS6ZJTJ7MR55IPCbpQvZSV1LQvzSSpXkk1DUO7Vx8TQGDRgQM
jP1s7kL2IWLpQtKhHx+sM9RGEJb/4rxDaKMK7oV5jo96U/YgZYsZgPSDluEcNGa0082iTUQOtiIf
DKuOBagQ5xM0+cSAZ6OmvX1AxmmGX2DkWEHeseBhKcn2IVbVjRnOEoRPVG5wjwVMzhMgwXzV/idg
6As7D6QyQNjJh4KDGrzPq254D5odgCcKnWPUT08pOY+Qka8DkJ24VJp8kaYld1Ikmf3kvaF5wjSn
ZpgOMS5Vfn/q0gS0O7mQRTOAGUYGhf2AiU66CSkYbQvkeiLkpKr6Dxa1MkZHkjXh+5Cpez6uvrFe
3Lb4y234a524JJ6iQDqJWpRTtZUvRXRTKJrt/ffV0kU8+U6IUL9Tzcm3kRQww6/Q0ttsjbMLzhXy
Wd9suppBN1G8YnEnPE69iHZJfHC9q0ZePu4HOILIVPjoMp7klhdlxWv66ACNCuX6mS2hujsP5EKZ
wk4bTi3Jja/CmJPwRHTrA1OeO/I007i1jLjkXI3vuDU/0p3t4wyTdKEHfpP0XGBjGm+gAYalblOR
jEUOOllN0zjxfyWMJ3WWcOMvba7gcwtBGXutu9/k10A0garWrYKzKoOdQYz2uTq7sQ9+TtBg/qkF
I67/B9pJ3AZX+uSIJJPr3KPc3p/nzuyiH03266nnq2qhc7bW7NtR0esGHnTA2wJ0vYskcnxL2yIL
4pxeAhONhlZZefKMOWQ4IMR2jW2ULbeVUv6pK276JFUiF6R2Tnnd7rJ+Ymr+DpLWVPNk1wtp5gMp
Re3tizZPyZzOd1pBERMbGu0wow046hWV/j9qjqXfc+bI4fIjEtIoYMoCOgdM5u+1/tzKuRHWolGE
WRHwj83ViEXsTD5uET0GolpXy0LcWHWGOLc8KIy3Kj6PCJ02uns5fsjBHmVSAWfEuf/GgPpzilFD
T6TOqGuTOKSrl3sXB7hkgXaWkhh5y6LPyfeqqb19HU1nGCFpi4eZCFJduUpPWIFeDHPpHXMpBvVl
+8RvtqHwAHnSAoVHL5PQ4fg6hWpoo8c34F1gGVSwhcHn8cmBLi8X9C8lp2L0ZsVHLeYPjiOjk6pz
Td6a2RToTbW06ScJAWnXvnnu4CEYXozW5exIyYbWb0qpzietJYpfk77mgHA+8RTv5A9Du4e4WbJY
ylylA5mBa2jHB4gMfnOL4lyVaZcvODZbhDexFNJlwS0nkylIJCQPzlbbZeiVRbwGxW+jHubAaWT8
Ezn8TIHQOb/vmEQIdkEESsHECavr7rBn6xCUD9sswr+mhODPrWEcNHapQRAw+EkcFsT5j0x8LG7A
FIT1rGXv9zl0kD8WdNImm2L8wD9fpveTnxomhTcBDaiZKybiANazHSetZlZWbcVWPO7gOVsFsHPJ
Z+OKOwk6+x8MlSS2zwBzn3smEPGbP19iJMJ9JSWmSQP6kyoc35bOlRZaUWFB6hLzg+DHoeysBb9n
4xCF/8h9JPoh/uF1cKosMV/H4V8OwVKvlWO5HkVOZ0/9ovB+o7rl0qpuU21Itr5NyAS1MjZj+C5+
llCWBnGlY2ynkvAzN3wqvFRXZL0X06zyw2r+wZVPHHMnR6H0ajlL4R6GjTugDBsKY0wULy3xtbgZ
i8inG3oGUv+bGaVVIUEIottgHjyYJl96AucwSNx6DG97R+xhVUwzMz3stGxRhnJb47C81+wwJ7nK
+eV0oWeFK98cAQBoR+oFjVp67mcAyUqf+8ecnqBAFsZmDFXgSIAqVgfbU2pcZIxF5E7wIlcA4yXg
3y262FMkVlFVeOYj2oxFngVmy694AX/FOLqqZbd+Ifc7torPV4tpH7MVTJ6Zl7NTiRLj0saWFLsI
l/ol2S8mOmlFGMiGoFXRuE7UeFJQZXnCf9jaEdh1ax0to/l+XAblGGo2gtGPq6QVZvceObtnJ5hA
3OeBMMiEADRv/D7gXFYkB8ki6HJctuzbaqIAajW5hP5AeRV725g2Me2ITZwy2Sy78V39jYxcfu6F
T19lyO6jpU8/Tn9onGedK77Pq5iolujgI+FmTuem3yxi1sTVCMEFTSKP2fEnjdBhx9XbfZbvdNZZ
2qVB6CaeHXO32dMmhFPlj9CC6DIAX8yZQDVItxS/mR7819RKrmgKnQKzJ91hAC3W1FGrwJvoKYJW
RlfcVIvTGhAkH0XcLlkhBGo02N3AtooXHCoXZugWjYDzL2EubFXbbghT47wnZWZr/15cNjmVzlY5
hOndNhZccFxmXz8Hhy94SboayvWkrdUlqLg+Cq7DKM/d0kvbeOxt86ByDVM2x9sPwMtuodRQFDUf
+5/sW+4ghM5t5p79p+6ATgLpKWxk48G2N4BYdjDyBM9/nWFnu5GU8EiBK19zbrNQTVvB4KB3wOTd
1I46YajlNb+wZmEB61ys41B2qVKQQIj+yt/Wiy1X7ndwQWRr/ptc32bAxrUdVVioGDJ5Gtxyryos
JHvflnTiHoKvwU6CQFCFxsnpQrKVT9lCijkYjymZvQu/6vXYNwVXye4NcO1o6KHvDMbXK5v7Ux7d
Cz7CtjRuOg1sZxYdjuoghJ3ioB8Fz1+58NmA0YBWU0acAaDXZuBBZNunooWgL7BbsOUDpyu9ZLRM
nGfWVNj0wKJOUur6pn1z8hsx0L1wvaeuxpL4+b0LH7dNiHFDyxWIQZgvHSQpAic7E3x02PMoKiDT
bX/EI52bAd02pazgksykUpbZAKONtSJElxgrHQhlx7i+6xgjDF0MnZoaXaxz8QLniE+bwNqGS3WY
CWwPHDsyU9/gKzA46B8pJ8YDca1WLBgWqyntcQEvsVjG3BFdI+pAq9934yeNZceTsQT4FbL6fg/V
zn4iokaa+ma7GbfAmws4+T6wgWAzpMdw3V/mUd92SoIUUAWPKquKFQB+99eZMA2UQ8ejfjtovf3/
CcgR1N92cCDDKeNShjMwJpKq419JzsT1F6rjK0fjrAiwVHZ32Z2knEpf4Z7ehqNKrZllq3gVKVzk
3TagpUcZX+V9ETYU9PiNHmAELYUjQ5G2HtvffiAA+4HV6rOn0CjIExr17f0+d39mtaO2YmgZJMvx
Q2f/2os1DdUywM4Xirkr7d671I2iAU5WPRbKsxWt07GjQBu42dyPHR/n/bISahCs2Pwmu6wElF3X
SHPsga0XcnjHOfNTpdyNg8PD+WVTvx1ohrXW1SI+4bQas+KsdS9WviLuJ6AmXdTRtpdphhFSe4UK
cMgkaUtxMPfo1p6rlNn0EuLbUDcqBthFD9L+09lMz6px+dIxbeDzMSttAojpiCLkzDf6NpM+RilA
nAtPsAPYvhCXW9D8wpTmLwl3iRXsPa1GIdy4PwutvudHFh7H4FkjSOWm1+SAii9AID1eZkQYKAnS
l2QiHao6h1NV4X5Crh2huz4xDNkLy04eTmiapc4JYdy8OHbZTeas9vGjo62LFYTKPpu9Ksw2Wv01
TOR2rHIkTRQDlqq2E1a8r5k0ybTap6DmUQN6YiHfTFTeqV6lWLMwIxxA+5EbDmAATaau+IxyYxs9
t1F88jW7ZbYsCGlVTXtXx/IR5y8YSuFUwd4ahgHV6GrSyao4dYARTN4QnvSY4dxS/jRPfAKpfbZH
mVTtmsaZmH7S+6gMKa6GuX1+w6Shs6co0SVFiBHXAN0Zp06YiEWWbPjFemNAozeoCkhvsThWgF2q
igf23+cbVt0DqMy+/AylGZIdcVOAFwHSSK5ktRKcCpDYdJ6dYsEJClXJ8Yo0HCc/t8SWAzs7/uKR
hoJUO7+wBTXuv11MXCFObCJq+okYHxFe7NIvTF3c/jO5Fia4rLxIxCRSiJgHkbl7qIHtdGia6jom
wyrLBxpdToaocuiEGQvjMqSaws1+F3hBmmfD+mqvOAUMZ0XD2iz54N6WVAUCmpYFEnXF5lhPpM7o
imaNofN5lmS35U9Es5ABgT48ljT/27bdmtJKtIahnFMFnfqTy23XTKr+BDGNQS5FJU1NluYaYKcu
sJdK/PKg2UoMRmKAoNpZRsgFh+K/2lyzE1e5O/s4ScCZCvX0IA+RzVm0MSBL+cE/K3kvNwvA172i
94AXW47vFKbsTvvtBzPCnRMIEuqd+e+Kl7NKPEI8D/Mu3v0Ahq1t+++2E69HKIQiLZS/pO56nrOS
Uup1865h/TcRPbS7ZaedG0eIjDmXOdQgA1FwZCvriGFCGFFXjO6ebV02bEfm2uBslJFpf5lwzjgo
OQGZfHyDU3qjDw8PUXFSL7/8C+RU5FxnnlXE9WAb62DhQe+nV9Sx9i8K8yM7hH4obZbyhGAsftRQ
zhP9Oa8okcJqzM03Yx4XtNBf0Lcw8Fo0zwroyJPPVDQhkq2Jaqkr2++Lmc9MZZHgILToBP5RqiZP
Odku7yltAPJbTNbbxFLPMi90H6LBaHS/GnmEl4vAUbO1iw1jvtATZG95nuSiQGZW8qV5cYsMoW65
fvxV0bttQ+1gfhnCSlInw4Q56CwjMF1gFya/id0oiTuWUuQi27SHsCcETUtUbwDg+kD+JRlRwX88
7tRJWlmmLHYFrK4y8dw3wMwn9E/JRlRoVGNhI4IQra5Q6fqvOzI1v/V39QkX0L80IcuPHO85OORv
BYsyIJzGtkNGJmExaf6uYndsexfzK9t6UIxiE1POvKp3ygdwqAvXhpR39rElMXMK07oX00MTI/KU
HhGYd+6hAm6CS1iOm3SPrXEnsgb8EFyfQPtpdykwdS4pqhnIqGeHINoR4l+9X1UXw1UFrFW6PeAw
l9aQCPqv8GArRny7U7isbncB3qq5WSmjKe7MerFzM1t3h66Xy10LSYLOw5J3hgxvqMs8Tu0Dcn12
MoXsscms5ALRgfZdcstcmX4Y3L/Rd0C972xpQjADvV/4UoU4LNkfVicgKXn0xxAZkDFgcjsmsO3h
n4LafFbXAD/ugDazZJ5qM8sBRsBVpiICLStG201NXLaLNzm33xkyczvnM84JHwbxL0m3c6wcIqAc
dOccJcqi5y2WyiY9cYVhYczFkgO2iE35J5RYi1FAtEtivciQAgMOHFHBqfK1lYVu8uDPmELn8MHT
CAHuDygUyI7Q2JxAd2ndJK0voXij2lEJ/hLwDDCx/TvwB6wG7sb4+bvJz6SbhFwSZlfFyNCOa3eX
Q2BZGvokG9YpBkDK8wp4RK77uFIv348qcyX70YThdZ4ysZHtqyKMFuA0AdVi0KazUo+Q9OxY6F3c
/0PCuMBt1b8WhFTf5CkME224wMOYd9vGX9MBCL/Gd6IbSl7LYy0WYyTbNAHVEZ76+5peF6tJ0h02
Qsth6DJg8NT6KKM+rR8kELCw0hc6FJUzJMgB4J17JeRipoYKCQTgYRMJA7SLADIilehbVD5FogZ8
wNrS6zEgohwhhiIOaRjfQ4HMz7Qbg4+4jyzu8Sr7ZL8q36500PGBXjyTQqu/LNiUE0ceh6UdLJU8
M9igd+5BO7LFAXcb+nxl1UEx8wlBn4NB4XCPkr8rh4DD6+mNHR7FkIIHFbXpNhbOtn2hWDTsUxQ2
r8uL9AADC6E1GoZAifD/6bkT8Pdt0EettEA+N+7/9TXpAeuwZnNoD3xofdaPtJLcPIPepDUgdRGf
cRhWtJAbLCdhvmLT4GlmEvTNupqtFi6U8XoFY9tTLsrCJ/ZKKVo8LTiX+hIxqaeaMKVAVMc95v3a
ya+rOGcn21ZKg5SKge1ojusE9vqJQzDiWG0IN8aJvbR411HggRqKzELzlHWRsLjWAMLcrBtsR6eD
4ZTSpThmWqtOgNM7ZCK8ZViqAsrwadResKRvFV2cm9L8Me1OGOxKikDmy06MV3q2UQ1BRgZNpH2P
m8GaHw6zIDPbQF3po8s1xlJP//YOoUnrD0FKOHgfYH6A3uCQfV8vPigfW2JzAIsG8vaWIzLKc7Ov
PptyEnkh/zGYzmz+/Dtt3nKuSI5bEmTSyQZakU38hw3xlbfrEWwLMiLkt+tjbMI6WwXa223jqng0
zwTw3TosMRQB+oY3oxybSWD5Yi3DrOIESXdV5VxAYGtyQpWsRMnR0wfSDqDUtNmHcKjqdHy67Mao
YwuHhOFL/rFWH1RBxwr/Utk1wUtToON19TWIEpI2u+bi2mEwo1+RvAER4SvDrSqGiTfhO5vQMTOV
qFhyt3akUpakDqm320kZcT6DP/SeWdvCnZapGLMWZfGO4bpdoWvtaXLA0seFgjnuXBOUbwGPK/OU
jMJcK9wFTMG6XiWeCxkDMYKacq382ZptQyMbNvFEZsPxJXoJMZ9Hg7b4BRsBQAM1t9oAihM18Muh
m+jt8UU/9i2SVjpleT0k+Y0QoDAssTqXOH97hOVR7CGN7WPgF3I5BNSqGkmZyKJn7owLyzt9rGtk
ewbTzEHn4LmYLX4F72JusAIZPZYtJ9YSpfkaIJw25qwE0kSj3YYOLgtXRrE51v/FU/seaW1lmThf
XTAKaxf9Ac46Y1tljHOwa97AMI3dDpDpcn/BREqRL17njS/XtXQTpX8NyOUB66/9cMpAYJtl26md
WF7Gz2V0OQ1YR8jmyOex12/6gCheA04Mum35vxnS0atk0VTEE8t/I432JSZF0HQqIgQqey2xuRMz
llus6jQCUa2cTzR+D7cBpaV1oO9P5QBUFcHKPXE/0nrby8omU0S7MAhHJqVHzEdWZrQ/swbr0CJZ
XkeNblc8AbBHGY7xSI/HNKvw80GcrlaSGJ9W1yW21fRFBl+iOBypc1JZAe1B2PZXcyMk+c+wQ5bm
lezqD7ZKxpmyzdOUBFbmRS7UK978r8Nq4lsvgUiVC8k1Ptb1zr5RCK7CneM/A3qkMjaOO2wCm0H5
eWAcxqKxgvoeVjP2TjY4E8enx/vE2SxcR8pPtH6ew/r12GEeDZhzIdsOWaY9+HXTGCPTUKDLGEi7
vc9i+W6N+Nn5Z8+P+F0XXn/wg40t0ixhyImPEYtvM7DEWe7c8X4Rw+Xay6Pa4VVVKbQHI9x7ghIu
k7V3RpHa+BaWtSBBpvAEaqK4zHG2ZsyHa5yC6bFJZ4SrcSXWXMg92G/Mote+r+X1GIIWoPvT9EMN
xrvQZrPuxJGLmzmhvmzKvU0Ww2pkpXse1/1O3CbbSj2xXJNiebZXk8SgVd0i+toZvDH+HQBmagKo
DCRYFlLwL93ZXVsmlsammIdy7jKUF6IxzcsiE6RVgaw93wrHbDYjooweIOKYYJQd3Tic17l8rkTv
XTXcWBfuasXoTsLHlpwf0jXuhcaHrhZv/avsx+A8jZyRdYjwvW4u49kcqWlislfaPr2EgHLi5G6M
n+6b77x07/52hNm0gzoqBz8aKmtkGMpkgIAbdQWZNH/QT5jklsgoEjHzaXZicSRZu8tzSSTSmAGd
LrEpiELvQYkyaTGajesjJvFLGuUSH4O6xZFn40ajYcJdC2B9WMXuQhMNCvTx58SBJJcx/5miiU6Q
qkjOIwn2fGAHLQrFRhcUopQSsh/1W3ILUkfa4Tud1enekXdbotxMwAMl+JHV9uLVkf2sgG//ihB/
PeAfi3ep0nhP15+lfd2OZijA5KEy1ttiz+WfOGMbi1bu9v2IorDnfxAEggFyRHF+qOi4bLAqqW36
b2hNQW5KNlwrxoj2MFxDPC4GnEDG+YYHEVwCO9IiuoU9z+dh56sgAmiu1XRHT+gCuz3/Mf7J343h
MHiOaQ/qxuaoQDDPbOtYd23C3qOv11Rxxg1IipYzi6gQKQHZX0Uy5NnTCIzQBTYfFjnj7Ty5T0dW
t4eJHpC8McrgvfjOTb5nnBnES2IIJA4/Lr+fC8AadRS8VLJEvq/nLXpkrlFC1zYgnb9lgXghaFe7
gYHTYOCdJGbQMuiWII8kf8YeICsvYE592l9Kx2VdvQhw/4p1WakD1sJ/kCgFTJXSEcNl3KT53KvV
DEx9xUrlm8dHiox259CZoEkY61BuDmyd6QgLUuDfZQt7TEevapJumPTavDHm/Az/GOdHpsVTDMiu
aFHCpLWwixu4O8IIn35yRkPOwR/K+iSAd1fVrKl7VcDGN0DDjpWpX0oXQD45kLSVQN6WLB3FAxSZ
ioFGH5s96LTomVCi2NxDGVQlf27omTK9PiMVHoh5vE7fdJVaRyilXxY9jZ6G0lvAx3yXp+Zq/yog
8A3u4SUJMYpJaYkZbZaepgz/LebkoIQmdu3SHdDuHI20xb9deLfxp/zmkahPpIs+O9cJ95IVV2Rf
VZYgjwWMxNAaYopnetcVbTsBF+ePm+Tu5DirIW82dwvncDSewP0gTb0ufEpTfmqyUOtKV2YCeDLW
BgN3l0ntR7424FzcG/oVxr1iaY+sJZZXQG6uRuq5uQmRtsqDwYbzw7eKLjwxSxnbX3iOsk6ZTmE9
y00XO+9HoC9ISf6WMWJYZ7NNdIMULDk4SrPHQ+bsaeD7IM+p3XF2zoVfsJjf6G4b6sGsdbp7GmTe
ieDWtiOSXPL7OrvB8+mNGwm2Yf1Gci2Ylg364bULtfgJuIHj3uVJsB1YjfhE7a7SKHylwDwZau23
naucqKfaCRl5iWlBgo8DSNqu+hQy3mVgyt9J0QpTWYclWsiFVKaYA/IrngAQsxyqb4Jful6oNaiQ
0UZmtUXpKUSDF8dtx1GAETWB5NjopoZHsBvlhLacnpPTnmYnOyQVaJRB1y+O9YHeOLeqk6Y5NuZL
hk29unX4hYlIqgWKcDXrA8oWhRRFRlFBaIY86Rx6OSF6IZQuz558C5FTo2U1Rvl52y9+UtuFDCQe
gGibrSTDV250Sv+Y6WbznYt74QP2pbphvkYxIY9M/8aYH1R10EBAEGp7T/SkYe3vV/1KsI5orZWe
omP9JlCPzJMw6hrYZDzkfUU1wdh4l6L7AxBDVfllJ6Ixoz6aZwRmwImGIG425ZjBdKeKt4Zx6895
nCHqww0DleBKzlPphhFk6EMK9X97DcNWiKRhy7SQqy9FLzFRQ0l8q5ct7N5aUR6/z5r6bPy9G5Ii
HexTzPhD21VGutaw0SccqZkqg3L0iRrHrTTE+VnKiPy455fvv0Ao8wXonnDfAPdXPkRkltl4RY46
0LI9TWlRTXZzPP6MP6VhA8aZJy8BcqHvIMLxYK+bIU2N1/zOkw14037VamLAcnW6eIxMWsqxVtvW
dwvq7qPkSfbuKiF9BszY7mT9ma2QkSJ05yBJMRF3qoUd6nDghQlQx2J/KkTqlCkSLvLTskcwWeQS
yreTSg9nNKZFsIeSgap1QQxIWBdiTBsnx6pH5dFilFE03R6nReC7xGnO70+lzjBb1JS1QdOWEJ6m
wtiwy6TF3t+3Oo5ff7P21PEr3vquFEh4GqqG6KAEnDM5OGwm2PMcL1G9IhzWAsr0Kx1R4GhV/w04
rYNlQ288t9xZn16oPXyN9azj1zKSDJqoaZXPeF9jSXKL/ThE4vfmLygzZufceAJXN1nVoSNLj5d1
XAzJVgD1N9ZNRDYIPN7U/5t8ktO5y6A60AmRgpH/W+dy7l/FK2K2meGPNasFYROgW8HBC9/YkmhI
2nopmWrAf5r1/9GwikfWt4JMmxr7oiNT7lXr4SuAAW2V3ObUbpUKQOIPHqqa7AUoF7d14PRLbhub
wUrAFp/J7q2AGydmgxh5CFYNFAUgaIozxlJeT/KmSPUUX6727sWl9ib0e8Td4seCjJJlSN2YMose
smqx2toRSUKRF1ctvpHhHqZVHg9ErE9pUczemksKKx0GOpvONft/3iiG+ciOhR6Mez+jaXItbzg/
VRAjzdFcnL7j94HuK7wL7p/ZMSqIpk68sYwjMtz/9tJzwp+DBo0hUrW/q9eTaBSIzDBLLmAALOEJ
JEERMdmYaY1SGKr5fccDdDlVrDAzZJHmHVhJCaupntfV2MdFflQrtqYcGMNlh0S8Brt6lQ7lu9ck
TjvcSvewZFhepoPlv54rHIjgz+bSiVJCe03HilsBMDAsqGKVOuiNm4qrJw6VjbGV2l8l8JPbl4Pm
HWzcaC9mcKSySV6qMbIBkZK48mj07DcJpPl3aLe24ZIvziRjPr/tasTP5trU+byQhZXTYtpM/ZH+
n0ogLcS832+8hNF3wC37assswXOqjseTBVTqzn2dm+hY7CjZCzQHvUxnGaopvCtkO6EiBFISX2ux
pp15MjuIGSX+rWlP2Z22AdBQVD/ojT2R+E6zsGQMSeKPa0TPBRXk9WQnfXs50ZZoBWfedMeA7P47
YBNYfiJvQgWWvN3U1g9RZOH7uNI/GXb98tFFW+zoKpRe8wYavyn57ccWBIS2Vn2w79DqqGWv4MZv
5hBHImIClo/sC0LyaLc5bPjGmguxzTlziNrRKSjoE0Zgftiwr55Q39DVmFjcA8gye5v4Cf+EvrVf
+YHuIteemkK30l2YVufVRQK926wV8RSoCKmxpyrAJ+YrCpZPIvpOMTToTUgEIwzysm7gmEAtK2nb
e8LeO3l9C7vcqni5fN5jl+4iLYpg4UnHNEO5p9SL8KL/2uXQAUljtDYjx+UfuVymfwZVgBnAOaEk
MoTElIHJ1VHUBRT+3Zfl4urT2+x9Nm4GYAn3iDkHsodcV0hBz+Hn/i2wyRUTplBhpJqhZ09g7fUm
rgituQVSfwnNWHUgAPJjSOWsH9uTO2Aeh7qxpA5q8MZR4vriFWDeEP3FO8xPuV6YFN/xd6PF81bA
LXnQC8uG87dJsuZ+0azXAKKF1KJoAjOJLtnLMLeSmZEs6i4eiP2fJItSS+BlL9iaO1uMBr9Ed1xw
X3ONDIDh0ptActUxV1AVSdkmChYqrsLnDmhX/tJ6xKywpGG3EsHw/5/JxOPuTFqIClMSyqxa1WoZ
aZodLmunyOA63WIRWuP9ve6XTuqK8jZjVLRgSqdWHW0YPZgqU1YA9kS3O9qZawKVRj3R/nEKviCH
W16yvCD4kgAHREJjNWi0wGtJ0niJGE8mrsZSojZ/CHJ8LW8ZuAm3yoGkdiu7mbafquSmwea3wVee
VsBZOWuYG10+ej75sJYBYw1EPTxlsNLldQfjFwFH48Nv8d+Pi/EQwLM55NNkVxSnaKw5pz2+0J9i
SHt7LMKFidyNtAniqNOvAdxChTmI59+OlZj+Bu6nXoa4gYkOLYpKGe7k7x1xO/o83kG8Fs8E6PVB
UDRno+3HzDBk746wywHx8JOrCjUzMQw+9OG4WLyuITIRtATmR5PW8EuCxOAXtTACm2eyc6UjRdis
N2yJKted2t5DHYwG2ECyOCmsRUPPrg2Ri32KKz223LA42/KiakiTbSR1rNEunI5u+BqeQAWZCo8a
pTHl+wB/O7ya2wSkm70oud1IDsRnHAjYpsNCzs2QZX+N/MLEr8g2chn+maydIJU58ylQJHDMkoY1
Kv/sFFYjc4QgKxUjuM3N5kVgW/yBwKtT+VI6PaLsmkQUWkKmCD+uy12s+R6MuAuSRpkukgrRgLdr
777l9Z39nx9xaV5is42DMfTwP1Ue7msGDTNwrQbo6byXA3E67E2ThNDv6h5uqyDYublSELta0n5T
FmdSTCc9op8MeMUpoFx9FUtMbUK2lLab9XNQ5msiSTTC7Z/BAJRWkj46P593kyoAEe/TPDS5vPcE
f7mKDb6lJ3Pq7/eDm+UQ6e7eYm8OqFuX3r0uXjAFrHY8zuM5F91RBJg0AilhVuBJsjZyVdxjJgtT
fI9mTPL7kZVFdLLganQhQHgR/i5VfYzwI6PypLtne2IdhGUaIdyISKZPJ9FNnWBloDAFnAJpb2dx
6kS+rP1qs632Uypb9PwG/ixRO1DczGMpPE9oBL2bpZSmFLZcnYkRDkX+Mtqte9UsywVHNR36nSr0
HX+5B7VFHVXkOaB+SwjVDJOH/jiPMQxYub/nB6SwwGGn3QIccpYFYUE8dnjz1jLmWQIP9L62HWC0
o/b7VzXtP1zReIf/WSubaj3KqMfxFPeRRfFZzepp+RrUfU5aqNVUitd5WPIP1JjvFUt5CYx9EtYq
RyeoTiR1GtTWXH3t4vBr8YUp011NpVK0w/3RjbpOWlwT82FB8iewUslK83lBIansiPpB8xw/Ay8H
K7toPf8DqBaxhKOtAlDGL/Pb3IqupP05Lx2l77fRYnP/s+2sprX5yhZn9M8vKsOwXdE8kjLnByLl
8+RGezbopX6D9tIwlbo60Y73HKSgvBMLX5n4Ei4kP0oDwQcY1bDnH/X4epRBIdkrCa78yHr/f70h
P0Jk+EIRA+CPeWLrWZ6o14vq6uCQS441KiahMlJXxjppIfOLnOnKBP4VExSYbX8LYhWuZpb1jf0h
XpyPV/k3Tyc7Euq1q4DtEhMVRvunGom2YOPB8qH0UOt6Hmjsfq/PwyJk9k9LUnv3iiQy+r+CBbhd
yCT4iLyBDjivo0C6rS3Ord//85PGIkX32z02pAHgQeGFUDpadQ5mbg40rCvww2Oq8VTXNSTQZNLF
yzfnXcvncGDG92VUWSpVHFNfgFhXVUJdZYfOIrzbENA+P74In7IDo+RyMUuhe7eVeGVVO0KhU0Sr
PZqV9MShYfRY9MsV2h44vIb7GwSH+XnD7wXcN8DeDRmfJ1MEIVU2rxm4QuJbPIhh7EUSrMiulkif
96foRkaSpUNfJaN4Awirr9zY37yZxH5l8qlvJSNLDhg7c0JkRa6EcaqMW8lR/bCLcG5jXHGnkUDL
nan8Uvn+Uj3r70An0L1R4qWjkh0W4kUAGw2IvA3aZw6OyfNJMfHgK1Hic0rjWOI4YtWvaVJJMaPq
lyP7oYygGFVMQJ32MaiUBkt7f1vN7lWGF6hj+cO3B9Zqzu2/FuMiD5zniIRRYXWv1Mx98TDDC/Zk
EIc6tzMFJXXaHz+0pjxoHtyVWYh5am0c65eK+55ebr1lWUz4Q+9Kd6ZQMLh/xzvLVp9DimJL1HPt
q5Otzm2NUtmHEsRfgpwwjh9m7Owwccv+7nEoqUy34szPnDPpKTVRGkUHvAU/LjyIcCq/r8zuiQTw
1F13qztaf7IB1XvYWQuPRoIXbfIUya7o9wK1e7rAOHZjtU1NfFgOuWBVeDRwNEcKb3swHb9MzX0B
KTI9K0XbvlIsZbpfj8expDB0ge9q/T4HWUk1oOaY+NrmwWSvNNaXY8fYzWPyDeQ5St36zH+RPePG
6nshkDHWpdvXF2Ra62qNX0N/fY0gZHfZdWmxYgvoiOn1hCG/b54BLS591eRGqurgwd2/Don8Fej8
EFIW3ICZ2lJ3Bz73KlbYTtxbjF87cIuDVZard0oYEsfZTapu5dJ4gCv4OZ5vbE1YPv/QIGu5iMrF
+Ti2lviluCro13LbcYaf3l5KPi9WmkTqJTpl6cNv16CR+SY9IhOHgYCKdqVfE4xR99P9gUq0Eo0C
2+42uo7mH55WKIQn8+DDdo5VGCwpQQ4Asx3ZananfhICYKWqP2ln1LtTilJhSKQka1l7+N6yrbHz
ySEmAPLKdZwIK7Fjqb+IFVYyMWz8uKitXAJUrZfo567x7OlAfLjRhGZvQrVmYcVH6m/EA2rA1Dgw
VXbfxuOcZC5Zd6cftaNt4Y3DpMYbZeCpuJpBOBaxXdSK0fv7tBfo3rVZtr8gT8kr2P+Ba6Gi5fdC
PKNioAXdteaPOiUVLyglQHiGb7l/dj6Ms2KtbtCDiJ1pr4tXkHNkNXy3fnj6Qj5UyDvwxHB//A/C
PEdxhcvEnGGwFfebJ8HNxKKHT6YKvZAEc9GxtSYuVgzpXNzirEvFDdRyQeg8v5W2HfwzxILC2evk
LSRb0lH/7PDS0xcPCaXhxAPgdlEVfjvesfbVzKv0qs6pjJ3KbqEtsH+io78gkNmf/t19uwKY/szA
YqEL4UJnewZOx0nz405DI5miN4DhVO4EA3Eo+E1yLwkJlS53G92CFzs+m835ZNS7poJzI5Fd4AGv
SAY/m92F1PTmym5w9bp2a0j+2j3GcyRmfGmIADFGdTCCMlKi75KU4ET52aZU15GF+thOiya1F2Tx
XiXyQ5JXKEXt19WlYJS3elvipD6qcB87SBHYX5doyhEMQG7IGLPSxN4JwkJ9aqVn3cwVFtQW266X
fvi5U5sCo/bUfsscnqINjrJigTtD/YjGZXa1m4hI8BseaC/Ruhhlo7O+YP3KdvO994w/HULI2IOO
SmHnjlkKUeer0aoD24pH7sW8lEcqQYz+xfGNpxCuCM2B4fgAHIHYY/2hZhNfUwjmP4jZ4hAM4L8B
dM89z9DaG38mxK4S9w3yXgskXftKQmTjtyOrH2ITPm2ybUyndNo1ilzOYO3uoIdUUM1UZajz8SUD
q3Jzy89lEn1c3fhfsocQWzRyrO96e+OpU4yxmKQvwuCvIpTA8ippcV+dlS6XGUQFZukRW+ASFML3
JsWW0rfIiPRX4X6TrDraH/s748GDoyPFcm63MXR0diUdvIDlfmrHWJqFPhZyt5IbMC9Knm75eqH+
Pl6eczacgeOTrmUvZMf0Upp5NbCaaR9zURS/1izMUWvwMiJPdS+BFIvIJvNCfrmaJa2I3rDL2nsp
aAmKYpAWNukQ0jq/6UNY47rWee1Dzcz+I2pX30e320YKwEDOJ3WZmUmkSxVILBG2h0lxrKYnwEwY
hAzY5nx1xwfGLB1aH7tjHkjlkfqSQxhKcg7NjlJVtjv4E4x0v1HxllUUYqFWoG4S1jMIAERQFaX6
UdsWLzCopitNkPlJNWUIes1gelJmFxsu9PgiH1uV3stdVOD0B14jy+klWL3ZaD3/zSe0spSfK8Wt
7bT2i/K14+5SZBLY5x/N+d/9BqNmCuWomZnZUxy1S+tEtLyXaZekF4bs6qVWqAo6FJTCXlFv3vpz
fLE1Cwrz2zNaoVShHNBK7VdyZQaozSmbAcMzCEkmc1xgnQ49NT3G/xaTmPdBBdoHj0nbOTmYO8e0
SJ5Rna+6r+GrsPc0Q2XHPXAucm5AZ/CE4gVMYDcyZsrSGRpS+R26ykF27ckbmGTpJXZ5i9p1wRzu
EGKYQpKYljuPcVW5T8C/3F5+rXw+C4wE4oYZ9tMpbRH0kBh3etHp95xDjeMGmcrOQLtLw67l+7iW
D+PuCmywH5fpbp5lbWEQyg56J/o4H/LHrB769+ffBshlWDcFZPUngEd+QjNzTVfOgBMFv0gMlrYG
5LHrZp1sY7v6voIcfty0EGICdb3UdBUCm1frx4dXXvBnESfPkravuAsIaZL+OXfPNQ3ZkGMMy255
ATvvBaweauoTfwASvC6PDObFcPooZSQCVCbrIqD1WpAjr6WywWQiahNxnhQj/pQhizlSDTyjlOfc
Pc/fbvaqvgSzrctoB8wZ4yHsrx4z72JPdXa2xwgB1yxxVIfYWQymQkzP9usvsl2bDCryd36NFG3L
xe6Ib8C6YX3FfeSD6gBqpkt32g8JUoXz2FXhXNK+djQ3cY8ODJ0Z+hnQvK3LWN1QERVmZzx8Bg3e
2lxfZ83KhZxK6zB9GRtMy6bsQ5cHDlgHRgAkdnbW3rXMxWgfpieV1d/xSENu1HvTj+RltizuMsgQ
S8UWGDXR989NQlJZZZSRSRgbUbpQZfQ0WHQtKAI7KLRQFY41CILXkPurSwTO6gvc9jbxi6xtVbmc
cPJkHvBA7g/gvlDtbGZcWeMpM0PR+sAITZQpqvlMCXZWzV/87cwIePgP0LJ7Jlt8QIWmIlMavh8H
U+wzGTNiFXdCXAjEPHwewMTPtnKLRD3Zq6WOkLX+ER8IID1yf7JZGBrou7kz37IDYS7iSUBufFfy
4SxiaiPKy1i5KlEyFRy0sBBkIvcqrow0NX4wHXyvN8WP0Ujcz9B6oa5+6vj0Y/hVQQWY6ErwV8qn
rKfsX8PRiYpXRgFP3U3fI/bkZxgNPSGMblC43oUiHsVZgVEeHkjTtjoHlqecE/ExZksM1r2ahv/a
aG5WzKFcN0WB5zlSENpIsNS725KFduo1rBc8zGVM0ab3Lue5E3M/3LvGyPUAZSYbhDpfHieSUcpr
GT/tTO6oIbJ0F/6MJPE+pnKPwDMJbQNxqzAsYV03d+o3aaM9vrPtYDGVQNoCQK0BFnbMAs7PbI5U
bo21VkizKws9ddkTZ00kw7LJ70RlrstKe6h0WKNJR3opK+aXfOaJUluR7/EMPXUwOtfH+SvWYce7
XQZkxgpGk6WXI3W/J4OfFuEuANHEIG5ObAOZDEMRZUOv55n8BnFs+eO8V39b0wqaBFPpeAOYTZ+W
LEyiDyJ4laZWYlc69d+SDwt12ZttmF9ovCbPHewu2OS9GJqE9sjK+61Zmy9FBPOA8mdqW3pVtfUx
uUAZCWQePgCQr/k32xtsqhRc2vMIAcj2ftlB8Di200Ub+7b6ryeVoPEKIsrtT6vcWmmG4Ri9I6cs
TzYn9jVFUvF69E5ICaAfaMulE1cRJyilZRCFuSSmfjLJnMOzYLqo/4w/jz+r2xV/HBFLuqP7V/Sc
nQq8jtv/QpolwP7W6sYFi4K2zBFzVtvlh0pRKt4aFoMONA9pRr/8DIWFb5hDKadyVBCmDTtM8akT
Sy7BH/1lrgpedzfCphusAFtaxvRlokvZVvIim7vRiA2YQXIphnWgkaW0X8Vf/aOi4rtfY/mzPt5W
t0GNkIP3rUEoEpnJtJpvsgUTQ6LSiwLeV0fOrcWeaJ+sJN5XZ5l1CLCBz8QeS8acnZTySI4SGBSd
+ofgZV8/Sw7Bmvkaag141Xbxe89ddvbkt7JJSWWlPbDwpFM4E5kIQntd545ypxLtlyGNTfyj/Iva
v/LGx44SFZrjWqbr0Z8ThDaje1xFDH8LfqvM6B3MvwKLu67IgK/KWnlypIMDq7Rsl8FGusp43Eka
FI0DO/UCMbTG9llOlKZ0Br+d4JV6+4SKiPoSuhQAK5dCIwTytdCSy4H4L/19fEHPrZ+gaRFLOa5h
Xec1bEbCU9vBNLStzAdxZJNrfFDiPSmwXzThtpWH44Oo8+DH3NBcHRP9eLMrtb6cbxhhBuUn6vH/
aBXhQTxqWFB5nlDAJ0w5Iiz4FajjyZjAmbGcchhHQag+Vht+VrBRBdPTcXjybeHBZhjf2WM89Csf
lIZdaEAmeXDaqYMV8KYwvEfMSz/51YlIPvYExY2hkxpV1zzB6JKmAw7bdhg1GQl9rA8QonSusJpg
nsc0U4gADSYphkpz0asHL/74nvxvO5+itDGdZb7KIoLcD0iluE2oDl/GlT21S0bx8ZgQ5BV/AKax
2uPDBeLXo/Llsf0tW7lKxhLA41QqoLqcp3VnKwvZifFOuHzIHvVp35lM3az8GILiMLF+7DTGfiRK
8zIuwha9E/pewMSJYcXvMTmxL5L4Q6skLvcUHklJc4G/Sp2fnoFK566+l8G82VDG8ZZTHapKTlgz
sZxrzQbzNns6Y0ymGfW6/RvltrNLxbn/xsOsvllhvN4VNVgv4Ud/xxf+iNy4+rJXV9K8xmjAUusQ
rclp8vz3No4ewdUk29/F9hNL7CoCN6eFVr0Jqukv2EidV8wrMfu4MgKBYFOOC79ajeodC4xzB5BN
wBLdAQhC1qFPxpdcAaFxu2Wt+nQMqqmq4gBhvUlrbQ+G/LR7EBPzxazmuuAwgljNeozt3fps7Hhs
THDAmQMYuVcTLMMr/HOKKiHfRrKbRCZjiO2sLvbxLTkVymy5wd/ApuIU0ZvhR/Q/Gq1dqP63MSQe
dTjRDKTHYJQJSjcdomnnya4gXaxsW6wzhm/pCWNa1mR8lXEyl6Dp/hKD/yvIXtj73gEtvayQ+Z+F
FLF3JYsTLL9BhRnD4a86RnMnIDaKaMm/mDF9BCnuHSibf5R1/AGlefZOyrWhIRmaP8T0lZePEAtd
7CsQF30YQVUBrJhNryJvFD4beXBz9LZZH1TMc29lxXfEd2qHrEw7Of0XYZXMpRQSIS2svPkxJSXK
2dEXwEeS+/podGOviLyaR3YA16olQzhZT5dlosgm5lJSE0H9jeUflzxLQU03SsdMsexChQdZbiOf
uf67d6AamFVRi19THPSgmYHxKBkPIZSYil0xmLDzChDlrUlWqWwcRgNekjxQWx1yLYoZbYKPzNI0
CwTX2w8udiaKTHFKrwS5dXF/DJVkY+scaHqPEu2EK5PQSPe8WUCLfggZvP8p50cncUlry5M0taT0
tMFw+LJrJNTrbTpeJiGGGcJfJeH42N8Nty9AzJYw9aO/N63CLzS0qOTyLqUQb6x+0DJqzY1w5f1q
32zzV/CiwTD8duR7d9OoR+p/wxQje5/z3jrFrkxmZqsVrOZlhT5ECZ0kcfnKRqSs0aTSD0b37ylf
B8lkefidkB0pMfah/wnIkKRC3Yl++k6KgpjHqVMWAIGAAiH2UHel57DU9FpXOz+SOlEAsRwkryFH
BA2yiIFgWuy4pW4h3i0h9AQLuI85+d7/2JpZurmVtTp8IfO297W+NOpynpd17rdA9rYyr5/G1QVR
76KQO/gB/Qi1I5F284vaGpKrhxPaSV8yUtGUp5HM9w58F5S+/2+mGd2r9EFSUpbp+eVP1v8mxOTH
IxIflViYNy0rzJd6N6XTR+m1aWzh7eCKZIg8m0dH5LTWpDUDbLHHSj2ca2NmfAuCTEjrfnYgfUkX
b0eY3nRYrmo4EZsljxSkCbEUsTvW5HxWMLoFl0Ezt6xHHdUjfYw6QX597RfgpAi8KVL8SF8/hSSo
MVXm/WpQ4ICF/n6R2DY7f7C/yiLnzBQTtZABrmCqkNM23lw7hD3qJY++6lqMYNy9g2EPegfzHbP7
Ks9KdmSwh7A4wVFRxvwLlGkR9xMOahKJVMktcFPaLdVQUG1GhwWUbAbm/LNdJuZj5y3f190g/BLQ
WzDge1JbFmj9YmZepvDpZ8HqYrFyGzEBgQWAsNsBfvuN4o/QVRanKHtIaGh0bT0o32RKhJ03MSaj
a97t7GwNYOBc3MvfsJRC4XTfLZHyave26m6sHO9fvYkKLFw/dCkapftCCn9AZaeNxvI0M/3+cJgT
FHc9QgoI9J6Fn3tEfi/38F/tNIBnnTIpUWiY+YveMC/hq+yqAX04OU+6+P1EGEzgd6xhS1Qrbwyh
sAKhyw9cDXAoGaVN2vHGLOZwuByD5jrroUo0j8D6TJ5SiYaK/kggE19xQJXWOxT2mXVICCC/lHOg
DQQwbpHLeg+GfeHZA+3xR6Ib+arrKc7dcOWfcKNdn13nmkSKfoUJmsxxah2z9kYxNqU2w/wEbo+U
OQZ0XmeenjuHpDARzokEOgnM6SRcZ+6FXrVG8vkO6joueScYQ6JRGL4CTi2Bb1eWWoPPk4oi1fgj
aIz6aCllOiBDDF+4Ma3IycqS59ce+aLidAYn8ehu/ERTGrWqik+mM+HHmHN4zYD+iUtBvsS6m7xq
CqIvRoTItl+5sMJKIaAW1vQWrEh9asXTU03E0mRbsEF3G9+INxgMp7XYhYrRoYFArMGmNyCxLJf1
5kVD6oxycFEAf83W7BDWutWQK/g1vOC+06p0k26kzYq1OtG1E7W4ecI9c1+0Y8uyz0bMXVEONcch
utikU3M1c49WAjd8rv8pUqvcqyvlzGcn3aNtyyooLubV5W6IYk75hh/12qVxZTj9ztO3hMIu2Ziu
ZijYH/7o/jeQwIGTcrZinNnJekEQQlp7JfCDEdKCtqj1rjwl9fhAauq2l2wp+x5O06UXeAZglKP7
eVhG87GHu79/u8jqrEQ5He+YcKb92kWTQp5tIATDLaHpFKxz4zn8OGiZocBbgt+qkgnTDS2Jn8cB
Wp2APK7Ew+FcFuTK5N2/Ga6rxoSl/DOSCbt9fX/3Txsg96/L/pC99V5MVhPkem4pquffqdwullS5
XC9qloMCLwnK0Bo0Qcn0B0L13kW6Nl0nBtW0gOZl1FaJyrET0gUlY67WUEDY8Vft/XVk99Pdveq4
eC4ea+AGaFyzGUIkJFEXuja94KcCy5GKmd6Tj6QADXJ7EeBkT2A5Q0vIp+XZ86BDQyvgWSKMVXhz
wcSDZLpF0uFWnF65/2RbBBWZV/o7DV9+jwy+o9pdHagx7rUyWrHKxYAhvA35dipPvSu3cP7BqReW
tE1SDrZb8PAVR02JLtH+vat4fJYZPtnjJ0DH88EuP4iadi3Fq77+x6P7nsdJK5BS4jSCQTk72XdP
Zs7GQjATnwRmnME8zSqWGCMaAq8JQTSI8Ni1spSk9lXeCkR4F/jpJbxXWOKN3LtMVSxirZVq5Qjx
AFjffypktpHhq0juwPG72CfoAardrsEn0VVL7sSZ18eps6qjqhQsInOQax69EM9d0VE+DVUtHzCL
jp12wIrQg+UzP9f+Cx3EHJaFfqYywvcYHnAqRQlzt7u16dcGJgLRDiRG3O0BoFPDEtgACKA8mNdw
welaeItRCKGjGv1/4eC42bEIkPyEy7K9tH//vUFAkmkHJTa5ntZJGEPuNiwFa6MFTB8SJnvCV1rU
aH45GHBUwuLXHTOQkIqFNgdNsuaXAwfZ5jEOUzYBvUSFpmBUG58v/QgOxKEZI0SNd68x83yQkVca
UsZfCQV9g7ocZQTrmapIPi+O+Ev4kNf8lNS9tHj2LG3raFm/oR/Ad2BBykKoeFiYTZBaNGD/gj+d
R7ol7An+IHTsOVIBLvZs6Vu8Tf3wvUffFKqLJQWiyr66aBmfaSGm448GfIqK7FasfPDDNr2AzBdD
gGFVYWyC1TgNDEP/LmKe9GObAH5qNHtuXwPP7nvbU2M0JTgzyeE9qj9pejBDFGtM0tDA8FtotxpR
Dqci9iUnhufOfGUC6nRXHl+3Pk7vPecTFQcwmuj6Zd6NsousMklFQuSSgu29CPbfrzAphBPrOtd5
4Z4PBVtAPmtYwjJv2fFrdleatWaPh7I+yMNKIv7/j+q1qG7XF8U+9xfEzgYY1YFwA2Qs6DT2UBwA
SvymxmBqexMnuwL9j45WSb9fpPlbhMwk9nlqXou6GdWJPp9Q2yyAONUbSsqhgK2QKqo2XnJYX+6x
2QyLf1wa6KD5X6WDi7YhsZgfuhvET3iB1knungrLSzBnv7sNCHNq08mSTESdS5TDk6dbZkRtDkLs
agam0C8g6nv5M4DAnS41HZxNoli21gOY15CI5fA4mMK+gL34DwaAMOzBtcEm/L1QvDI1YhfEyHiZ
+uQ6ipmvOToPpt+terScyd9kbzIt3OPRGnofpH7zQeNUqwJcsgPwoOSB36R/VQqI+kQv/Tc+bV/Y
BNrP50v0ZnUu9L4mHa9F7BSwzIylDDyvXb0qoG2HQnpVrYCwCsRBc6cxpesXo5kJMj1ilddcmtMv
Gf/h3HVksvwj8hxsUDJ+VwBEfNJ0Y/iVwxFHipuLHc4oqTl8bRg6MUW3WiNKp/uzCLlIgbR8MKEe
GoDRPqslS1wtNBhyBiCSkoQ79kaOIcOqyHgb9hhvnNKpp5oVjG073JuL53tWP1T8zRqh3jvdLl8U
78Jm3DqbtesJhc+Jnl2dE0+aRJqw5Wgxb7MdjRQ7II+fDzS/Mf3FWA25sK5nZihwtnUru1inK0EP
hVPmv+qNvpzY2CL4t06hhYiGmDStfBffeBbDKVZ2c4h9gC6zMG644bW2XiLl+cvT4zixbnqG320B
CcRvqhVv43HueSjPM2DUFoEcbWmLIetPyBJKao9Ppu7gZswCx2DiOn0pByQaDXFFZHMAIuyw2doP
kqo20abIOLZkp/6xFwWCpwJrEOctShBtysGUjfzJjmpDEigta24kTr+yuQwgEJjl2SFT7C3BIDqA
5WEs06l7siGOzjWBlJpyyDNR1lyXn3GQlrW0X5exap3eREVbc7TK7CZipkpyOtgX06FktYx96RM5
o6WEZUoKxrNqiBrhCXYegNtqBoqK6FFJmxiARvWPonxvH91bWV47ZTfUwh6VCFyx/+pdOvwnhw42
hjwUvcHfXfdp/394+QyxQ6oTT9ZnS1i0hrOFOE8Iw8p0xGcqjfA0ElN2l2j13WWsCM/if8jt+tBy
RFGhX8wjW+anCXoD8c/AWghS049NLOhLqPGIB3/HkIAT1WNuY/BwAlNGKjZ4QE4cOegU/vXO6OFm
FrmN9IEBOT8C/dJwQShje5BVwv0scNINh1YLkHWzpJiykx8h9HP3cx+jMZAtkeWah86iPSkit+gQ
NYrH5ADI38ajyZyNugAQkeFneWYJPSEyknUNgIMxImYday7TRnqQ6oQf8ZfHJC4R5roFJAPV0g2T
j0I4bO4y3Iymad045igNETIqbIdZb+4OKSUpobWJell9/mVUyWluhvIn3faMFBYWXM28HtYvm0JF
PfD2Qyqx7znPOVJA81SlA8z5WEjsdz94lfxFZMT1OkFpLRLh7L658SR80WeSAfReHoWI+i6PBsoi
1o9xyzRpxiGZNJnYFQfLk8YvCtrJEuAMiFqc0e8bsWn7SX/zFlmyAx7OHFhx9ls1XqjKVusy11YJ
lzeOUsLsrGNnKgpvOUo3HZd7ByjA0xJmRavUC7Ma8mqWWVUGqKHhTSdxoXCIyD6DDKjlWXBIG19k
kGPLa9dxg+k3QOqdMwt4ll0KgP65yjS5uxHTG8KJ2Bl2OciWxPH4TAh1KRDUk/DXOHS0JwyXS7Rp
T4xoyKBdFjtXjC0mOPYjQBZ5gkeWQrfQCby6X5f7MZzx+IHH5qGO/hT6aWNeNMn3/9CquuR24dYk
gDldpQZyK3h0eSyYpyu2xPG0z17xDI/q8efDuTTfVwtBdNy4bTNmq4/kVRQQc15UmUloewGfOGHL
YUOgKAHZIbwg2hrGNj+3oHfkOlPyujY3U+SGWMDzbDA7wId0QxdTEr9b2NeGuNR3XEnfS5Ael/TC
w6NoHBmsgb3qJJXUgFqMOxOlPbZYUN8cpwOoVME/s7mT3VvEskdoQ+HfNkAVOcqM6UlMSCeDFn5e
9N4NEJnADvR8qnrYUzxz8q4oCFQsXyrj9WebRdY0sWXPVE+NYFV8wbp13ZslXLWmuaBrccQqsjxi
R5EA3gTFic1HyvPrGkK2RuITpIWoLuFU61P6B/fd3sPQ5KRXJOl3GDfFoE1Ivgy0FdDh++2C/hHN
BTshPkWmpCpvoGigDUsIvvfRBy4xVd47ru15hplMyiFnh+2rvM4DExDilqj1a82Sabr1+2qa2nCl
PldFJwxeTa/GQIeLPCAhiMqAUOEUtMBiZd/TaeXiUssSnWJTFbLX3IY1+6ETWPeVspeOsLi1FUxH
3bzRsTpOMtNc761ZNPiN+S1QiJACD4GEMPPUf577o9EUY7pVBmI3h1C8GDZFJDZoy74bM5crt/oC
Okpq+Bee15fqMgW2c+M4jhwD+iB+hAOjOFH2XmfEdT597AW+IEou8aBQ6pZtQWcRUK6V7EnnbBhP
psjsLgesOlIpHPQ6pTS6eWD9zMwVr/fgw6JpKfRmRdTeOMwfBZ92hNO/eDSKkCf15wxX9B0LoHWm
J2xDAdljtjmn8ZVc7e4Ldcu9SQMKIY+izkzXwM0kv4SqVleaAeHHNQ8CCiy3Z7c5pxQmNiDF1Neh
+XfW91lyQ3cR6xI38nmP2NWaxIFFOKeXXltQKrxBjGG0WcYpFDYjVgbPIoUxagg1z0qwaRBMZSiJ
oJaRQT4SFP7VnEOjHGDOtZzeHq2mKskJugo1H6Z4VmQ+RHDxMlr22gBrNg2fduvHQ5yHA4AbRMQg
M4WS3iwnqeO1/dreVyd02nUo6CbnEr+DdtpemaIin2BvfLTHCNP/uNXnps3+E+14qSgXEljJKYLp
6WdCLnl5mlrTgJyCSqz71PbosEGCjoYAbdQ1aAQNYLfW/aAU8l7Fu1G5VSO0fRZ7CCzmhXtFAgxE
i5gIYZi+YsSsHcrK3G+XDXylxTJe8t77qpj1FAVUh1v9rij+sSNzkWgicPS3FzC6sqBKyFlo1iKj
mD5mKUzDWelmTal+h87coK5aoGsgzKep+sNGlo4vPyVuSdo4pNx/1Aiv66qjjLcyuuaA8FXiIxih
EnT5HaE90b+h8BsJyPw/1e2Nkh/uzEe9eMbfkjW8ka4r7QMKqA2kRvq0F4+e9f6TAzriR8ImR1tO
vOgXEhwZ3ja1yn8vL1/Fo1QstmIS7E26HITw7pqbAUDdGrUlPYSNM1K5fFlDqUXpBmzSOAFWNFcC
ITDemzkD+Uypg5qEGBPA3Y9rAah4BIrou9QgEVpzjx2W+LZ03cvV9qobN2wmP1TSmNmX2FF6tLTH
uJrgGA/9hXm6yEMUdxVg/HvKky2atffK99j0Y4TTJd4u7a198bczLdhPNbjUqi01/vx5Hhxft4AO
00CSqpHyqpQNZah+L+YzRjT3zWZrfId9xxnTxEnFQpMt401h522VqvFcDAvX/9G1XUNqkZPaAgVt
pQn/Avrf1kuDQEkYoH4ly8nQJD9ZdqnUXehMXZAhhc7dB5ZVqYLyJ5BjskR24OCGBbgVuzuw/z5m
vsI2wJRoLVhkOAGRY/0d/nVd+dDfpkOSTJOx9JNQ9VgDh4Bb01iNbLSrQ+hju4eZOa2KGSli+Cqa
BantLU3ru8T8jAthSe4+1GfEVf8MRgkqqG1XfqMEVfVO2eWEeyNF3QKQZx0Vukw/Ef/DGI0Ozfsa
PePTwd56u+awqTsF0uhZgYF35vKjNn7WhpnMdl7CX5WxnDWeNebwKRF7kfeRNW6K9VRfxS/06GG6
RrActQ1lvVv4rDa7m55SNhtF0bcMMGK1mVw0ELrLC2V4/H8RIRyY/tUYjvVjzSLft6qJsCNS/yhB
BTmhLwviojxOBGoO5p/hdFQbYp5u3zltEb+C0o5oX3S6+uVFLqONdKw7w/hRMHi9FQ6mG91u2rRS
Z+IpDiIB9S7IPK7bcNk9Z/QzwzKopp8TEI9hWyBVBsgp+3H/n1vqJ55aWC15NWJf2HKg/nqAhwAH
84FSCQrfzkc60x0PrSc8kc/zno3J+ShT6WHvYXM6K82SekQQ/lOBRgDT+PCbhaMseqJWPQdBZRev
SSPsQmESVjgLZG4mjAmUfv7I7pFOYUdqOCuku1vW63RZg/oulRlvXve0w4ugPiAeaboIXB+SchHm
hetYczZuR9a9l3b0op79TNSxIUJiZy5clHuS8UjU3dgEfIwaWrZ42itF7qSxj+207bX7DCU8gCUH
qmcC4ypfh8NhyP8VBHinmxbZw8wCVrpoYasEfJ4BMq1nPIpF7kXzLbPA04s5IpbhkfUh5ze9G3eV
1zqQStJ1SJZYhhbxQi3K33V2AeFfyVBbN9EwJB4Gv8GgW3m4CYaQyshXibH41nDZHmCooDuaSxJC
JaomrimNU6dTvAjehi/o6u84rrk9UPoZwJyfko8+qh21XLVUs+VYOFc+TX9yysM6HhbPCJ/VMpNR
Sdq5yW3AesDuQK3tEZKUJt0JvRpJqF166KC9Zitrb23tkE85MdtM6XlS4YmVNZErkFShnAnCqmFG
liZ7Iri+6pbKRkeHrf44OtXstSA0+/faSfiWp/jTlkcdUz3w3vvye93CCvOoOVO94FnoeAUa+HlE
nVvAkg8QO/CG0aeRmy4sZGQ1FTAHL5zUGBDmrkXlVPPM9Rr3XapcAEv/btxLGTn+HmnSI2FLFhoe
+32mPKn26w3OmCIjwIV63QeDnvRvibZKGEat0APU5K5LQH6BwRzG7IWuNrRkDeZyAVKZpUk8Jhvt
vWWFoGp5ZbmKTVCAeyfKRkEw8qbzLq7pNopCNDqxk0HsaeOZFY+GcUCKJ6HTjPCfO4SB1ukdBm/5
0SB/N4DIDilfDloHYi/29ruVZ0f5LxL4dI04ph5LkVMCnMUN/YKt+8o3H79yRx1/O+BnSX04mjIE
jnF7x/rneggiDWkFAFjU8XP2yE1FZGn2JXwnxzRXCzOh4IrMermKR9kuOLkfcqogentDOkx1j1hU
516iSUO4MvAw97lDhfworH0SOzy5hvQ+PnZBFoGwdXszfDaZq0rkwqJOB4IG0PmbaU74F4+ISifT
FIuPb+JpDfORbemM318IfN1FnMo4V77gJcq/+ZRmowXwSYNkFiRoNTnY+wgrzrsOuORKHEJ2s6wn
YQU4Y+4cm3Ng+Dp+OSfTnjjChatt2Ve9fhCbCzp5OCEwq2nxUbgABpZugMdMZ6SgJ0XHmAIEirxR
ka3PyRc99hLImW13XlcoOJqTfELgCF0iu9q0vt0IT8VthSkqrhRJ4gQdPLQzucCscS/OH2omXkI6
F599ZRxszcQFn0p5ZBRBxUzRv/TGpRC3hZpCBr4ITncjLF8LNtdDDS05bLKWWHbnWbGQgSsqdvsY
XdCsv4csiYubZGDJBYyTOJv86Px8X/235J9YMK+wa9Pb6TEYfwmbn1dJu8ET2S4/AAv/U9IlCUXe
Jg6QWIUr9VlwluUlYNF1W3dkXFr6QHzXKvA6KEFn8AvAQb/l1UD9xKPoqf55Wv+0GotYVLOdgrlb
MnW6m0zgHClAzu5RrcjkwrHSRgxosNEo0ctuKW31csfBZme1V+mS0gnuztXmexvLKis8b4qVtE3B
Flc1DCINUa9sfOjRsTL+0mp+VvTZ6tu1GuP8+uBFYof17JKdZSUK1MkL8pb1v/Di8t3kmDcjFmtG
Q8bZ/BVuA0YOwcmNl0gfzOtV4AXWt4G1cLTc3rT1Eec65kRPrPo0uApHFY7nxgT6TRS160mlRwPF
hRGHHHw3QLD7mitylRlXS9RLsYWvNXHD0EHWrNOXXK69F+sze1+GCgodMX6EGp+soxnapitlMw3+
VC2axQJuMZ9D5VH2x7uVEmyaLO29rgstxVsmV8RU037WRet4cz7Qj0m1cBSJF1sGiT9el1zKIs8N
3ZQqmFPu7u5WG3DBpxvgqThoNi1ENhFUPtmq9Sk9vqXNunhpZld/YoIwXQxU4lytqMH7ZVSE+7AG
wJD9KTy2a3cVSN/SJ87VNzkQzoXqE8B8ux3wmochlXmIAnrbTmFds+ZjnteaYDmgP92GEabQE8WH
EbUjHQFZJuR7QmvvQzsHq0DX9cAkaI6Fne30LAbzeXOOFDRucKPH4HuuX9u4Wpiin22mSQ5zELYL
+i/wTekN2AFF4zBOxDNdhl9Y3IC2o593mGI0zIqyFFtAk9vAFwEBeDtQCmQ7wGv/QXbMT+deTCEN
SkMN0s3Q8xlAKolgYcSlmBqxX578jZuIzf6VCxYlS1DOTTi5c8/6UI2HAoJ/hOyPx0CIBqqRL1Rw
5JV6Ccept8kUh2qZMucDBwz4BRjvKYVaqwmWCIosrlEu20QdaDh9gY77pvJUoUb2IHG0s3eGNGrP
3L44qHI3XAct7+zCNpj0zIQIbXJd/L1DNFyaYDD3VrW49x4nxhmf9Wr/HfQQgn/686QTKeCv5zIR
senHf3WLD+8OS2pYJ7rUTbuPfkZv6U1+S57yMjAZdAo5lYdf87OUI28r0izzznZS6u/UqBRgKey9
uKw2UW2l6LvlTh/Zkl15sIQgfogHsj02rUx0eSY6dqlL+3fDJTGz/mMKVLlndgmXDwsM+ZyNsJTi
Eui4aN33o3ANvL+tVUEpVgVqhqIbMZQ3ITd7XbK2xW5usbs3XAU+/WkwndeWqcOeFsHBDPsVN3YL
9pfG7t83Ce4tgIWRZIJTe96SXlSSS7FFGUp0jr8NTGZjGFjTLCuB+WQN7G8PJixx3S2uP/32Rdbf
k/EL9RKkIOk3sLMbsl/w9qdla+brAd6GFJc4s6K1xmBTBhuuXj8VurkK0TLHMOcOaJ/qahWNuQRo
AGxjhd7oEqc5jO28xeMVC2/kR+GI+drKRM6RmO0XiFiN3c/DSGpbIDMjmppFlrgops+cA0q4cXxr
ythl8VQYaAVwImxzeI9J975mBGG4c5V10VaZx/1Okmz2xNB/R0qlz/BngDI4uNe99jleRa7Y+HnR
/SE1AhmU1ZRbDG0+yKCimc88ylGJledfwZe4ArEl3c+WI0g4/IaI7FSWY1Afffz6LXe9hmmCf9xy
K9XeKSM0Q0IlxE8toDZb6lWYGv8OLQJHmKMQoQo8WpZRlMCdBK+Vx6svDDlcgSREEuoRFla+AOEf
a+dczLHGFRhzxlHp+tAqX1RqduiBuotFt2EjBXCIKi/mBZOpi6NbDt3ud8fFtnHxrUpsYeNncNOH
YPA4Pm/D72yzCI+PV0h5UvYixTsWF+o92fkGtPcN/CWt/8Hfd0fg3uCIQUS7yP0FsSvqAJVw9ZY4
rl39KUYUbaUJpDR/M+HRd2z5dmyaVkUAwZnOe7oYvJw9tXg/7W4ve+HYY3XcHy4q/1hWtJbDKGCt
ed4MV6eaVXwb/xuqpjQT48qLqTojfgbXdQb/WViw/19/1+pO6tCLu65lc25QScCHPy930dvUhxI+
V0nSCUOmSBdtJ/q3zbBS6XP1/xZ9kXN6WZlYCl91sJWSR+hdJ6fJnBtYR9gRNxrdxw/5Gau4YXrf
FOb7lQnyNyAqSr0YXImmHboUru8tNq3WOFRvrHXAlaTtjMMY1xv0Tju6hZYEBghtsSgV+4wTLgIg
b+OuLjE4j9eK3ejhJv5Ab5FFlPdhQFyEYVWolhUmZmgcEIZoHNdauY+B6do5+8cQXT5jFR7M7g3J
w4wpcL3opONqCdNG4VYUT2uik/vCcHSglupV8xh+4C0I2swmoBanRpyj+kFTG/S9F19b3pbU6Ibj
AUmJbhJyuroOumot1IP7Mdad0nxPZetOCx298XD7DKlXt8wECtWAdq6cKX2DwV9XhF3FdFYBrbC3
RGw4GhAGLm70wrHV3bO246BbjmGqsfDU510PNwcGfhPNFfLmHkWKBcuZkEnE7Mq1iuZj+s5PmYOJ
ddF1r5qvCNUlXmXK4PSeKO/l7X2e965DV/FyJ/spqnlBDdRQaYPmbn62Wp2QaEaMXM4V2law1Y3/
g/Th0ZVlOyKsoCgUFkBZys5WgR/3qtSic0Z5hZK+kjIxbOkKUFEdzm1AJRuUB8i7ZzC7pll2mkUO
4ghu1j/9Zj+PMtswF49X6iZ+7OQtSiprHCN3pCYE3ssqeRIAxaHepRNsH+CyezpgBYEJsVG6KztU
Of8hzOW4IoE0GoSkaHbSMxxic/X72vRExAfebGzu7qmzRkcB0gecS0IJBqXvaNPgeF0xqiHflsOp
NLB9f+f0S+jijE8t2q4JnjGmbQ7h++MxJHmqydiKSsxY5EWN+RYoGyXmgUveScZwOlJ9ZLXcWLLl
dV4dYMNXxyzwITF5nr7wJWvf+OB+cxQH2e0WC+ooybBdoQgaLKmlVHRaBiEoFaezx0lE4gF2Tsif
GaU3/cBj0tejMuU9EDHp1HMZIzEfG2pijZoonqqKG97acct1tz1S3ZacRMd8KnBiY9pkJJyyTPTN
q8wMx6p7KmVpgVq5xcHu0K1SY6nCVBszev6HkYlMT9X6oGronSeETml+83KmCiXrTpcyrbfWM+He
jEYgGMnW2yjrP06ovhfSXNbyBrftG4OR+BQq3u/G1imbJ4bQTv7pXAEjGzI/GG5MfqzQq3kw35EF
DGdwk0hmqZuOiTsTXika+i9+pZ3fpHBRD0EAUJEAdM0S8PHWtKIHnfiMD2YBP8MGg3HyM4KHBnp2
JosJcBnH4PXVq+plLpX67Z/g/hTYo/6d0WEEiiJxd+Zgyefmo8zwujfFHdAKKgpF74ywI2FCjpRz
/niqdSGoeaPmEVzMsaJfSn5XBqj4ZXDunI3MWt6/6d7iXqx4x/LENeSzoAvU/CfgoQ9rSUE4O64P
ZHdfNzjRyZeN2SjX8OAfC0BKUZWvMNnRCMM0tk3TvhS4fUff0nRCn/8UwOX6U7oUc7lFcQcV7vfB
1hL7S5C7VH0SIj2jl/eScRXTPyNuSx8cEOZrA1VMIrDqqn3xAvlyLQhgZBTDp3yE8F4qADEVKG7q
AgeEtMx8HiHnQsmnClFZnwXEhvZqjiPODG1P6Zwx3RN206Y8hVab3FhmxSwBTs3s92Lhvhos1zrZ
kSw/JC0whbY1ntugVdAbX+yh09pqBAlhJWlzeHxE7cl9bcOtPkKRz8hlA8Lf4Ee3U32LdJnEqPV+
SWfd0SYpv3IrG61jNBI9LVEup7pyq7RtyC3ibGCpscUXlW0bEk9dRm/z0zUYN21YD4bX4Yf5BZq7
QpXCc1z19puHf+70mrU8tH0s+50L9RJyXRcHF5GrRExF/gx5wYxXaFMwE9DCXr5zc0kDlU9cX6iU
HyysDeMTKt902vOpFFSPrWY+iFRB65g+NIGhQiUMdE/T92AgYQx1uqW8G2NJpm5Khghp0xlsx99A
oH962pEHNSQWIK/OAQJsvTArO1d9dYHSllvsid0Raq9imYXPJgjnF7A4xKZBEwHH/97HWtIlBnD2
hJuipD+DHTGaUiPFI9TIzbAun4OSBTOF3NvKiqzgu960iRLnDj6parR5vB6Ml/Y9VJLvPlcZJbaW
vtmk9rCsQuAS/JQY7lo6s2bJzAYgGbqq06XN27VbtwLdCCZ2XBCgmd6U+Tb7M/vbiiMuZ9jpr6RM
mXF/x75JwK5RGlWbFWjHySOsgvHEMtyVt3Dud1U7MroA3cmf1X/+vuQ8kgoJQKO8DKrl/CZqe/PO
P9ZPHajtxchv5jTzlDSRNy1aMvjjO4Zhqw8fI1+IvDcavd89m0OSZrZ0sWeRY5o5O1YCkRk9yqXf
u0T+scmGz+C4BSEBhwP8ggEP+iNGJgo5Wl8aVo9BczUnQeh5fhti9Q+AJULGAIkiX0JtCktF2PAT
DYXVJZPL2/GHNmQjQ1GqqZtZZRk27hh9n48g3PDOA65zTq6BCNBSlGyRkGXvLit96e8Z8gtYSApN
MxAP8wzLMfuujXTsJAZQmtjdSmgrX4tlNtGfPvwddZQxmMD5eMQIJEnANg0wBWmj2scvRwFdR5i9
sd99GR25O6n2B1WbBc8uqEsVF2PwzXlSeq3xsZv4pGe4ozcgIDsMAJgF2nL7FjvO+p1ZIC646x/x
4IF/9gl9OlukZuNbVvii5vMEIHRgkbYxwnetxkPMlSN+TS7bSqyobzScSXRYbrRdcBpUlag5dds2
7CcTjUvwWM1leTR680r1q31RQxfUsF1ZNWyATIWZuOumUN07w5WY+75wi2gQJrdowKDbnIZWXg3k
MLGV17C9bG9tGqkdqVcODSGS77CMLO00Mrm2ulDCFKSniUPWeS2KUvpm9yWTG8rrcWv+3MMoNIcs
aDG2rC6GW77+hdRvt3jtqzjfbh5xKfousKcMxWrb/VkHoCXSB+stLwP1ObHikrhh7hCRXxV3/yVO
KiYJYkAJ7w3KnO+J8r4SGC+Cgki1TlW49fBSlFXMaCaUwFJB9JnRayqX7XyLzndpycRaASteBjNF
nTqjDmkBCEekSPpiAiRpxjxIjTFDAmQGLsgdBPET4TwCExDU7cyTq2ozthS1dQI3/MNgNe6tuS1z
8TOsoyaOsXFbhCPSEA5M1aqzJtARoiEEY6CVxNrgDQIMxukLHnOvrPwq+y+gSv5zAX33+m6XiHeS
gGBzfS2fGbnzJNMWcaGKuCciJIxwvV8dFFuj3/Q3hG1RT/ktYeRmSYEwDUM61C+mVnCjje7LGPe4
R570RuTOzMljfU72CB1QhOsoi24d07JowcRMXqtnVxW9yT7DLnFITw+/ooyku3XB0KLdMaWNlDqc
MIVFYcxloU4hL8twp6JqZbcB5IANGAyOdOiB/j+ecz2wz2lEnkBzQAC6ecJW3eHq6tzB9zyImvQ1
8EtNLsllTGX6YSeFoQtPz03PTrQrpbzS4MACeaX78mjXn3p43ZSWkKbBwBVMZalsSbr/haByHdZf
cYH9XIits+gYycFTlHvOMvDLaeEPu5rxspWJiT/OoyFCuNvuDjEV2MEYKShkBxhPmQ/y3b34fSnM
yI2JcXx0FNV+U79H3oaT1OaMiO9PMdQ7sdSOZVtdqH2nEGzXqI+g9GqQcpdYrl5y85eHlWBUFqlo
Wa7JcOy1qd3wtxax4JLdx1l6vAJlvhCMODEgU2vjDRYUsue108YzFKNghdogP6duQxC244UGm8UC
K6NTklpcW8gPtWSkeubOOEuOafJyj+QbnmOG/McVJhzIMeUVz/GJ1Kx8XMI1sin4h2hnZL6OKB/f
zT5mdGrovgRZ0oseqRmNgG7aTUb8EKSrcN3WNRuqgSb+hb53lOhe3bNDJRjr0yf8JYgmglBmZ/gv
tTBd6cVABaVkOk4UsDMPiB12E3VD7Bclr03D7n25AZqiavSVsCecL1xoHhq/1BDVjkaHGxRqk+2n
FLJ0deTQKA/x1vxlXMrAD7heQd9xHDHGN6XqUvdZ7Pa1dAir37X0pVbay5jbfB9zOFDpGQMcaBoa
PC/IWvhwkUFiqsOlV7e5i8kcFNezCnl/DIPIOEL33pq9FdqfXqwfdyMjx3mqHlBvdMp3b/6XJQ35
TJn9JzRBrSBZlZQEj0S6UL55vyO6Ut8JtEV3g0pQKh1zY9Eyx3Vrj2uuJD/4uNpj8sFFEPyGR49E
hfA7MboKeGTfvbafkJ8MvzixhXe5cuU5h2ZXQDczWhbkDyom+chX+OuJhACGPpEDLxwUCAHvKLwx
YdXTyMdzObB26mELHoEsLKeC7k/f6GbVdjz1HZHFyTEy+4A0MaMwOL5s3gQh/IV85ezbyXawf0vw
yZKhEtDQXSTWp4vi3sj2nviB5P6+qJDGkGGG3MRWpT1wXa8OS1TIBRZwsfd9JVTKgQhPq8PyIKOB
NDG+2rFl/B+xDhfGf7Nmo3F6/OmxCKgXVN2ocPPgrpKZOsphQlWOeo9FqOFa8+SP3FH03+3qJ/3f
d1fZ13zDn0TkwvA1VGhjgWHuKA0DkI0xYLYjpItULU2J/lBRukM/Ch1zVRsh1jwmln+ORCTXG+bX
VFE7ooLvQ8DXqD2LqKfFG/bZP3tAsjFLP2wSbMw2L35c3CRdthsZhmuHrULEF6aERZb1oqMCgJyb
nFVtb2huOqBPkRYvQq6z8gI2yM561XIPK8bXWWwutxDY8joTAHZlCl7zJDa8Mu4+z2XO/w3b4YAO
xPIcMqC2/0c9vViqojt5ZBLh97caIRFMMoRcenHAjLv0wBcOMbqyf/XQK5VGhXNvCFtxGMenU2EA
RqNl6qfz3tcAM4ADR67+g+nRwj68waFMRLWXrr54ebyCRYxGjnEFRmvN19iOA8S5p/KcxhEOURpl
k/eY0Wfso4o53t9mXw6pFwZ/AUuE2QUXayfLMMcPX+atdGWaVPfQtX/TwESdUeyAC8Ikb2fNJXVt
PlldYnrK6AsfDkcFCvWRFaCCFxEZeFhk9miMrmhPXHRJzML0SNjlVNLPdNTueMR3T/KK4mnTn57S
bv9wk3LCvEghOMbZgdVTULs2berw6QlaafOSvzsNeRkMtQyA9jjccHgFM/YrQ4eyapxpqsZjSYxR
JzmENKytxLAYeksiBqhMxPZTlvCnzNGyU+8VuTVL6CkIkThp9s8cl6XOLA97FbNR2PrBmjtWB1B2
7FwXuKvIMKCIcT7hDCOyqcgOV/D1RSyIysOcPVrZwmjmyhqO/ZzL8JAkN3+QizdunUu4x/ZmC+Ho
b6yDeufyPd3l4jFXW/ZV3qXtfoyayP4wz2f5wwSBFMv7joQJEcqtyeGHvorQfJBirpFEqFu2Qe8v
S9uJ1cb1U60P3MFZ+PtuESNFy1BLkD4gOQQrLWknwJ30/irNhZOy2e7HZjV7Rzvr48D5zvGGtxSR
qYSelDrNYn/Oi0IH4r94ChsgGfAjHJ3D6ZGFD6WQqmQNReGFfbWfGMHrT2kjQj/5jEsJvRpN5FQT
7B58SQbPOAtPskURTpnDoN4VurDbffZUaW+nNt2CkKbt+erSgz6174xZDxGKoYxMsQRZ327QOwDC
eHO2MQk1jhqoOePJV5acnDBa3Fovekc4vfely8Ty0Uu5fbCieB84wipI3OOv97vmFW/HhleBnAM7
H3zQLkNnBXpqHvHdr7MYOEpnfRbj2HfCzw9bR0iGk/Le6NUiltHvKECRU/ATMytWiMrZbHTtusbF
kT9mRkpfJknDK8MImF/M8dYhjJ2A/LDtA/PS45kt0xVbNiggo3fvaQF7P1MQ5Mci8RhqnQSFv3fy
96xS55yBVN3MM+a4AOIGB1ZJpTRZZ2eusG+Zj6StbyIv3aZVoECEUF2T4szt10o3ehAuDa1pEb5J
QkSGQ/nSFcXLtP0M5Vk6yR8d5kIa4pFxysm+rOuXCn07zVKf7J9OGegMaFJrW8Bd+LcDGYrT5a2g
s8UjmKj6gCqgjplDtQdQ5arIgHhDKphoLOjIukkXtzO48h1gq5fdZ0NeeNAyDkcYsG9QzltRnWnA
XyMESFMt+sST2PE7MPLdDOqZPHbdpatxhHJOUiJeWXT0jEVitlq11ufAnUv5TwuwDqVDVK3nd5Cv
u6uyJzX9EcnYF0hul2EPb15JVHGn7sOF6OxCr+ehnzK4NRdK623H3tJHj/Mg/wCb7w4vuP2auGhA
RvdbkYMapK4cI8YTk/gA0o+qPP3FSyem3h0nDtreU5ccU4F+auLsAS/+KObO0f2EU2/urevHrNMg
xWXETOr8vqkF2+kv+ymAW9T8R09wbzqwqO3w4TbBaCbzeJAAeINfYoiESBmLDS+YQl1YG0fkUidy
P3M9T9Y9AjlkFfA2GMhTVIqqsVsRk8tHxl/LPIEVVVsWN5pq3rmHsd9ShqFeE/uckml4ZMXb3nPK
/NxiRu5x2u5fBSES96l+wucCrlIEEv88jPG82GWfSovWu5XGTOw0TYP4iP+1d4gJ7qg/zPeLrFh/
E8VkSfidYeHNzfcpXYwOGLrHDxDWqt+4iQltv3PcnBymYW5XUTYRtc9voC2268SDwRZdx02yvYm2
ZtiZqF1PBRDTqdMKRUZ1TIAhsbUqkZSWqSSgxNBRsdo0bTYYrQSCMoCfhqsk0gXUE6Q6e9DT6BkG
bsveq4motmNwJhz+wDAVdWRr6tqOa8RCmkFXpLC0RREUIsOHvEApUyKPj27qyF3Xnq/bl1qmal9T
K0EUjeivDdzg+peZ1Fzjuo+eLx70SAB8DxBy6ia0nnru0FNQU0Pr0lfjq2YuCsQ9BlY0x9NVAhRz
LH5uMMl5Fdrs4mJJkWQwpIGw9QfUFUbGLmOtktn9HR77JzJBSesnKvTfQPSM+ukfzk5SiTnDDcHs
tEApD812O3TfnXCWX5+F4WKHcVy6VDlqf+mhVgLSEgB07fjM8idAZs165ztojUkhnULlPsaPfmqG
eF5fIxQmM4SlWfz3fCiP4sOpksxPtuMiE24w7067A12rFJw+/8XFy2UjKFaLIs6/eKIKcVOKX0qe
y1K3rtutGjVGGFVUe+t1MJjRfGIRSyiwezqFGaWCvUL5FmgK+IrfOoVYY5+Sg0Co6Dj1XLbYi1xP
oe3X14YcRd47NTxeQheA2N31UyvryFGK0zQVwVbc8eLVF+6MiOgXNMfp1bzI2TWlg6h5jbgl2iHP
DqlFPhztoP37YfKf4ao0WjH45C6AqeokM4EuPMLPW0ODjNzc4wqjOIW9kmY+ljLr9EC1RxlXxvCb
IJQ2L9KJdq8Ef9EMC77DVsSu0ZgIcF1f6I/Y1PNkhapcJJH6LaSu5qgUkKv0zmoBx3FxVRZpf81w
oQ02wg5miH4tcwv+5DnLGp6Ls6QL0zREMS9LitmByqR3O3pSdFgB4RReA+08ZTsVwwNQ9UYv0nax
5F4dkr+c1Ya+Rs6iyab0+ZWkk3KoFPR8YfaL4SdkhhJhxR92WXXLkpGGmhm91uHs7a+FMFw7OJDD
rfnUj0Pd1Roev/Xvr4x0yidiSIjVDtGJHL60p97YGAY1J4fMjbIF5T56EuLCZucg31e1yPDolIa8
ov4XChKPFRDb1HV66POK+qKtosq8/pnFYmidKkMpgegHmH+jkSibupNWEwKm0TYTN//Fw5A3QJ5D
kiSvELTeWlSQkRnLlMSVjLS/4lTHa2gBwzA1dI10ksqObVJxY/8vfq1DhoAvrFHInNOolqjF7hgs
FwMGNQsB7I3995rypfPtvxONhrnFGc3se/0+pmeYNUtbf73F78pCERCdZO+FsnBOA2PhKCwiWAm5
wQRd0foj+kxxxHWPE74Hg6YdLq9C6lsZgn5dMlum652EJIqnwA0E0V7UbEMf01akG04FB/X7aLHy
kFCiqH2RTarFVCBjwJQ4Jv1UHmqXTGBCRjCI/F5ZCEAX4CBX+7Ov3/pTzR+PbQsGukjIjLWk5pF2
2IIlWyRf8ruhzzTJsgKua13eAbXmeeaYX08E1/8sJhiiAmc/OvjUf8cKIDZj7WtOooaJlnoTX3kI
0HDeoqD0knNK9/huV5d8JuywJEn4Q5ABdy6E+455a/LDHY5Nzyidei6YpHm6GqC23eA91C39A1No
9L/P4/RKJoMIhQ6AnOtVBlghynlJpXwYRMwPiBhNIhKHYRLQK35RDVxf08QtGE0O2G9G1nQsh+y3
vINRhMFV0JQDKTm8ovN2G/vj7ypwHhEcgbsQFACcxLPgjneRZwQomkrLLjUAgdcxOuDaHJkOnPRa
qI0nc0gRTI233d+y6ErK2qpnHFpG4/b9sKCQLcsdoOaP1sohhEx/zlzdBK9APOF3l+/tnHieGnKU
uxgnEmWlmAp5PA8Xu54hFd+nUpzfdNw49yOfwTTM1Nq4gOfxISFs8Zvs9jB4iM+ZBuWRWT+3aDaF
HoEBCHhNM/LnCmVc7CyLSS/D1SRyYELO8P94A+QXDHw5XRnXpYp7wDxSpZNIilrA8j2OZeESunYl
qNMkJ4yiwmqDlEOcSoY2WYR/hmA9Qy6nZgKXq6Lta6v+K2c1vtB+MnBZZfL9F1s1ujBEUei95u7E
Tgmc9Cwi4HvVq8qhuy7pgIX/fex9RDgz73PlaNPKtu8EgQEjfUlWDopcSONW1XQMcttuAVYbBCNw
xRcPVdZQnTFpaWmqaJyUig/1qc5Y5YgorWpCxyeaz1WicqwrzdgUuQYQNM7kGfdSTls9jO6pgsR6
5jmifFsrR6WK8P2hjC+BdL7EiN+Mh0H7XtXR9F7CnyZIGWJbdLTtu4rLbgOfC/Pe86DJzgFg2zZv
S8OW2k7iQVSBSL+m5h/S3dPsPRZ3OP11g1DwNZRoA+xWN/sAOs0ZWqnr0QsBFIandn5H7d4Jv4M1
jNnhfm37b4nE6A94+PRuwG/7k/4xnHexzcmA5EvRGdYGXihJAuf7Soj1Jn3rhBS+oAiPvkGsEn+0
8uOr1GrF/Aiswh/VXJNAIU1EmlE/i4+qgRSL4okz0ZOOlTG/4TFK5qEHUqgIpSbJ4Fk14W7Vn3sD
x5e5J3nJZa36NRvgYdLoej7OKzOpLMe7rfW78ZphrhLEzR5pEERIlrblRntE1YfkguRX1O9v/n1k
LeT2RgnWNloI8q3tohXfCLhsh2yA8PcW0h4u1PaUqtEE+u6Yt0jWNQ18/6LCx67a0GRzOfQGlXXa
AFwMhUdHAFobLVH4oCLyEv9eD5bvnxaVByw1kvLdHGeQNuzOMtBff7TlawJEagru7KmXwPnovJat
xCRbFFl03x531sMJsJyr7Mc8an9Hl+gwMaheSvJCTYPh8Y+v21tH1sqja50eNM/WHZ4Sex3eunHC
xPyXM3a1BYWKutpVPJpGHlBhdIA+KUioUV2hWgi9ym8OtVwSsaXsotHncsqTpNJNk7bFEEBd/EYK
VGc0k2cueNCU2OG/nJjkHKI1dXS4aR+R9x17d7HFI//0axjq68meo9v0H3HjO5DIYf86pb3RgZk2
cDJXEhZB5ttwZlRarBwY7rmHaJDg6ci6mlRC/UF6bFhsDruvFXBAO2aH0pKQC/aSYzHyrbgUFpi5
O6BcNiN/rbSoEp8MM2FgGlkthXqzeoJjN9JcbMTPMQzBCCzafxbwy3S1Yzn5qhi4qPUk2UIHqujR
aYGEru6UhrzFUBWZAINihziQUrdRt0BU+bdYsx+WaEB7ZWESD+VxNozgbTqp1TmIaUYH2J3bniUJ
DRUSNUY3LPMxkFpQqodne6nzaOkgW/kvQQGysF2YYmzGE1+m4QKyxTjX7gHie6khD0Jev+ZjneVn
VOQ+e1ILvUrKW8j+WqD4pB8qNYjI+Wr/tRsSt8fToRTD3nIbb5ea0dv+KLgFUA7XHlcF8V5SruEa
m92qS4Cogld53V6Ouo14aP64VglkXMyCeEERul4G70ccaeJMv+iv31JQqe2A5+tN4pyrLYm+I5AC
JSJRyyEH4MA9ZN1Nci2L5AEFX+2OezWQYSzwH42Mjm06QP1FkW198cAilCJ0t5a/naapqckP0XPJ
U2bOR0ZIJEBTd/VVCnm0gprvAfC/8+U3acW5qTERanSZsJiFVmrFXkq8JWbt1W7jMiDwW03zTyea
QWwjedF3tfQLfib6VKSlnzh31OShEHPM2vbO5SpQagcIIJiUchYlXFN7siy6sLTLmg5jK2IPju5+
36qRvFJN2TVfC6O57KNiR6tgZwG5+1mnmcTK1e9Qmh6AZnugTbQncPKNXDjd3sQfOYRhiDrhpR5/
5ohoUOXEOubF/mfYdjH6Xhk2a8OtglKPB/dMIcOAGzCFtufcjrf9gjFc+wnytqavt3WsMPksuO+k
5ZIf4fP505+i27FHi9yZEcnHhDpwK3MM+F9DMUpx16jhxeeb1uObt/IUDuDyci1EhOlw0cI1uT3B
0yWsZd5ElRzSZ03uOylQ4lHe2vU0GixocE/iAiIBX7oHGfapsZ3jI3evyfF0aQBpF/MKHxPtTCQz
AebnFV0O6PJAdie0y6VENeRcGB9ffJ885e+TRFItblnLtm7FzaKYPSR+ieRMnA0+fo0RapDaSsFB
9TRDqomxS2izq22TtC5Zl91MXyxJQLu/bbWNviM8ZlgS8Qswgw/WMzrMzy9apOxFksJJ5XVoWrXM
BuUxj0SvE//tgRbfsfDSm8lOZBoDjZBGtpLMTRNEc5aN+JgmO8nZEWMlUlGZTRvGQgrGxHqK1sxA
+dxLHx15sUwhKH9sKceupEk4VK9EkZfHsLsRTMPUYlQ/CPxx9ud/BWhehsDO8/XQknY4No6yAQDX
FEMY3UJYTnPw6DDwrA9C09JLuH7KiHjuux0eDhkTNRO3fHdP999BP7kPj7o6qXKsq6gNkdH6WHGg
/tjR6XfCp4Gftbplcp8MOInUT8lmSUU1Jb3lVUOMcJ6YMiTKulMt8va5oGJp/W2HxJbx/3Z/KoLT
2TbadwfKxTM+0MoxaCPMNAi/AlyWdgWXzAv0Y0wnwXbfyFckan+WAR/3WHV8nc0eAZQy3gwr+5A4
0mZ33cUV9Id/qlh6w5BuZfpFginupGClk9wBpn9hgqTGH1oJdwWdPk1m8KyPTD4f/IFhLlsvV581
/La6zU+uKgKYrJIciJf6/kU3QZKyW64LbIm+wcNPouZrKP7wXXPQrHqRseXjJqJaOj5VB+QXLp76
S0IYXJwkEJdbkGs/ZyYEk/yEn+xJ1tiGc/g4Qj56ADiE8JWM6SB1Kk7m7jpDPW2m1dxklhV0HoJk
84QGAPRudhCoW1vVc/+0xZ5khLrBc6jnfVdSWYvb73YjsZCwfo6O9BAJR0cf6WPrMwtE6Ql6eAQ4
h/qieJXITSGbQ+Mu0sZbSkrC3+0zTXshq1Gq9SrnQCcxhnk3wGLhMW/T/YVElyZyNfT3uD6Y1Xbv
jAd3byBLw8AhPUq4jChpqs7bIXBmNl/Mm8jJEvAHpqlcUlS6RHAUwQEGk1AmMq+9PdSGKRIpdzJm
nz8QHgMC24n98Cs96f3VMotg92GjX4hQcM0ARZv9IBfptlN7FWQnuLJo4/zEYEbT8Ex57RQPS9ft
wWJx/jDmxMEGtTqmcVYEK/qlKHRuPQCPeYBMVwRPUX8F4ijEgScXJ9Jrmg+9zS8upY2I11Yxmwim
B2TdScKwVrWYDou+pKarSFICuyUOMnTllQxcJSG0PmE4biU3mXNJyvDuLeN4LjCiWxvIQ0AhX+FI
VefASx1LJRPAb9CIz1wkwqsENFc+k5ZYlBraBk3ViHGjfl3Ughhrlai3WVS0hcMgCGCMEeye6dzb
pP1zR4I+mT4hf7coNAKF3hTGrZ8hG7hNG4Ex29Afjq0Ck9k72rRG7l7OUtsYGsqrI8wqux1MGyrT
uRaCsLYJH1APdu765wqiZWJuHqgstW+n07AUZt8Qfnt+IXddamepH94rY4MCrfAzf38ApXGBzW10
1vZreLLp0sQE53/mw9N39UnGjgCL4qKibTaK2Bc4a5bJmc3Xl+2qmuCZNMixy8+nz0geBLguK6KV
ms+dAUAEbyIauq1SDF04stgROLS56kXhX0EdUTTUoq5uo3sc7iqN93zy+UGLGdg6hSZSPZe+yYLv
hPv+ytY8YBwcfl6huUosk7cluWNgZc1Jn0JuR3nvp6IWE8pHwqQpELJnfFFZHvABA5EmBhA0SjYt
3B8PUOWGG9EnpN/HghClzJJDGETk7fu1rRkkS3gdoO9CwL2BJO7oJvZJETFggRFTxtSWm2Vl1Z53
S1oIlmbyVRgUuv37TeV1WQAcfIaPYWWrbmGwNEjQRDUV3OE71gUC6V46mwcAEvJ50R/mgX9qoMRI
SKPbpgcZK3M2MQnXE8HLmlogDxx90D/msG7yUsT6HT6VKiQGPwBvY/1il8AvZOkfi+k9Fdcyns9Z
uUKuwkNaJbTyx7DrvQ5Mzd62dy5T4FJ1Lj4kfgmJroV97X4vrcjtfB3GJGrE/DYUK+Rc59tGTE4T
TWECR2+CuxR+GEeWmL7zou8AHvljn9xWxKNuPvXb1YYBanommAbahK6q6Id3p/BRseEe0PalZM4+
jzqFi/OiStUREKurJRn4EpTqe7X+pj33WjeV8X3eTtM96Z2YII5g35XbrgDEWcnTkCyM5SpDJ4vJ
pWYQwNDMGZVSsqBjz4x0l1lP9PXRMSyB2pX9xS8fyRpXUj3mpcU2uXGd4qxCYJp9XtyfGnxJ79nH
LQcBLVQEv/2dzb6WnaDB2YHzoJfS6bSPBV5n5ezH7G5Vn7NoXxzGi3cYV5SWsMLfnOgPLjg1c1ev
DyvZHH3JgYFdwRH50jYvAcPF+uYX7SXF9F3HVmGb+RYxQ3ghAh7gBUrCIT+gq7XGCtWfh5L8pnrA
67lUlsmGcrbeygmwFQTxR+h5a9keCsF652w5DGKv+2OrWkSDw6nGIO3V1m2QNe3fQJdxoXnNmK/u
K0ZEUTVoTKylzCZsx4Q7WRI9vJxrj7R4S7LOc/Af9iROcDqJFmSo6LFrzc8p/My18azE9MNGMrrj
VIJzPqoEloD2dI5LyI1lgnCdGUx6TPv8d+FJ8w2yx6WP1K9NZHUAYAWpfPAQcnGBIdRvyrn57mwV
DgUfOiYDLsfPgCKyC3bPa5XXJbiFHUbhV9l2EtEt5qA5wkKM9SojFcTMOXg/fekFmB+dDylZLmGz
sPav/oQ3yjYR3VAqHz/7wj0/n+JuG1Ho2OEZ3B1wuCSrCCWrPro+Si8GZScxQCQiL+gftpLlOPt7
iLuWbtZo8pu+kY61CulArkIV2hZS9HItBKI839VTPvdtojASICDDlRwa/KPNaVimW7o0GS0T1NCZ
NZOnVb0wonNsFH9TKWPAW6pp4QuWzMCSP2QHpyomOOSWxrzdFqQkOTBCgNG22nkt3YGEeLuCsXj3
FzNni8FgXMxwYDjuQ2R4ObGqf2SfbYPG92FdOGS2L9zPrVL53ynYAKxf7c/qlvukGNJ752MMP4Xk
OH+PWH7dp+9vS7VHjDRREAsOsq9BnfK20fQ/H9a+vjdGmYX3khnUE6F0jTA0J1uOVPcEFjdywc0+
/QJZRCKQAU5T7nJFINSRIwpuvdoXPGR58d/ydYfw1huij3B9Iju4PvcZNvERxDFUXO0kvsvJEi3f
BFVn1V7O6mZh4jH42Y41GQjaCW3mLbD07w1+faedorEe43MRD+jjgNJDTrUdujQl0bZ/Hf0QDmuk
7rFjYM57/MpClQnCwNBruqmxP75jb5NFRjDRmNvGZrh2QY5W6uGz2cOGVw19IpBai4+xHSJ861M2
IIF9W20hJJ3DqLaSwzCBqsKRlqCS0wN2wnOTff+JT4j9kRgwUDfsfE3uHRAqa6GSMxWQKdq9KRri
QbfitnRU6EsrYUplUFxW4BItuhLRiIBn3Avah+FnYJe4uzt72vJ+MjlSOC6LB4LvQju2ywr3zHdo
gXqu+/H9xLyveaRqxpxBkDghPybX0pXeLxvlq4GBuMkgLDa7AmoJiEb4E/u3hKwdjWxYbW8Up5mU
lKy7c2nFp1sigfOLMn8UIwFGQvAWcUhstA1iSdVKEgk4HaFm7OkYuVKAAhCo1u0VRQ4slR6Q9H69
AsvppfqIH0V+cYwDdv3usJi7UuRKVXryrpxyaPl8HrcJJFmvl0s7ARmYc0Bpi9x7M8UVZGfEH7sx
PEplzDj4f7Gr1j+kP1E9QWJ5DOcA3C7PfM0YVjCJEAlgNwEEPOyeO8UUOuqaql2F+AwjJTrX29BA
dFYwLOhPJJCRedMzPblw3xkC4vYKOTTAq90I8AWZNVVngQWShUF3brs3+PS2v1EpLm59xqd8Kcxy
RplC4Sesv452bbKS5RhHw/7XbS9natEf0x/dTEHxctkd8xHDi5jusmYa9y+yIyTsq0rigbDRBLMX
Xa/YtEMmS+72EY9lJqSH0oj3GEECeqORROUf4ggag+a+Vy3cCwLGSN0r/OMREZVeGH9wuGVZTzju
sopYFZuDgC4vsgYkg05IezpvKoShkggMC5TUaVHVcGOn8BKT1jkHGMq1nPvpZWID2C925EkB80Du
BaYZHJ0gfjNsBvHlHITvVEMSnSqw5gwzYzePRaIdqssH0vwvlBI63Gtf3E5X/HQ0suV/4vw1Kyl+
tkeCK8iJ63JDHQHd+qE0JFk2OKf36MKrFZBZVYap+EsJpsDE3m1lkGjsYAt6iICY7Q+71lw+MwgE
DMCR16ucIJxnj+ym+orrIMmjnNmeuL24jC1SkczDwgR44wO939lOK3MGQ/rruDPOyn7gTSyU4kaX
gyNsZfqvwxt4kfOLSghWdxxrIK94HdhNP676tpRWZ2vxjOsRqwFb4H3tulKEUjC4QKayMnZ3dJlD
XuwCpoNYx7o3iv9y5LIWRd0imxGc6GgnCc14yClS9+NDYmt47x0og7e9dkfjyS6yXUdJC9Yu34e/
KVKZuy6ge/fMhNWmP6mYYKcGxag0/sPT9N/ExeNwUs4fawJiM9IBo5AnLH4zf36DBZ0kLpVDhMTt
ImvGdkkpKVI8eC7JTzEEsE9An/GOhxp3pB7N/LbmttmXw0Y4kxX3vaTqJvcIQ9E1adZ7K2wXrnVL
qs847853d+SqHG+e0OPZ0JQzV5MQyOQxsXFQmM4PD33p3uTQ9sMbaz4OxSzIsGbKF1EnqDxX9NHB
8Eo7uL3//wH0Ds+8sSsJfnqEoU2dfsiUlBLSQa7I1GZvWSmOzXCgRizrOhX+/v2c090o0KZTAowM
oYVw1GaEW7rClwe5F14Y9CcoQFvVKl5E5ahVyqklB4EebtpMMa76AjjnstdXABVzvOEug3djU5Es
svDwa6h63RZyit7ASBvZKIiog9+symNB1HQL7TtX+A4BrDWotGtFbB3E7ZwDtJ/U34CT+Tkyn4/m
rrQiGzaOiG/w0LWr/Dd+0PIlDyYJsgwrkvASv5nQcbrms/18yOTMCgcO+l0c1A1LoqWWwnjqFZqU
1h3whbyXQxdOEJ53lrNtirDmoDb4A0N0Y5jp4Bzp6JP7IrqHi//Akm0F7wQzpwwWJrbbAtp9dpdf
yfQsQYk59zwoKUszOwYQvIKkSONydjpLAgtudeY+xNwHuS1qEEberPnUmYSnOUwq3p+jSdM2h6qm
0UXyaHNNzOWf5LnTuCswR8UKJNXxwhv4ZLpmW83bWxyI/+PQ8IpHxwdZVh+G4oU4YBedG1mYjJ1J
m25/a29DAP8v4mqWVsC4zf2s8FceMIs4ndWpzUgXxjC8au94PBIgvzlJ1m9rg6Z9PR9RVxqe0GRE
V4b3EHHVknKgy5TejmmMJ/m5BVKR75t3oQ5TGAE7o5D1S511QIl8b5Ez4IxYGWakhlqyI6Uve7t5
HkClqmbobKEkdRSC1lcM9Ph+BB+mCJssA6uuFpng/62TK08kgSNKBWlYG4jvY11LThuHoQcUGBZv
wV67Ua+kBMM7+wLgVmJZWMQZIsBnM0eE9aoqBsCY3/NZEqH510WviZu71CBCRKjlw4YazjJ/6OMA
i3Ypj8VPjZMYI7pSWoyzMyIGcuxbBQKv7NZfdsmRNrWKXQ4mkIWB8m6FR0HWP6OgLriB+37T628w
/AmLfh59ydpf2iCii7AHgRpfojWNXEr7k6rGA6Xkn4/YgMyOEXWh4ycK6vNRuZZkPJ6Cp/I2mJr6
7e/eidkc0uTh41Pg0HRY6smzlCN9CLOXsUv+aysAdjGvUX0gq2ew/Xcg8wQN1b0bOzLFT8yC4fqL
77kz06odh4Rr6NvTzbRVG/zFC3QIaHxoWmYOaRhX6L0UEC3zevkDGRf9SXnR3ljDHguUsh64iM+E
xnsH06qNWg5RVQsAkx5jZEF6bI/TaGoOkR8ehWq7SmrmdRbhK9MBlwhtAFyNh5GMX58jxEU+ytqv
yGFPdM8vEcf3tU3pkYcTfTAsmRkR87Q4k75sxsFUm5fGnhjl5nnLpW9JbfuJB0WP4+3FbafsFlvB
j0DCE/jxQsaL+GcRimLmwQ0EztxCRLztnz+0a6tXGZalO4BEuvobuLHXefZIfCC5kZULgRC+6NzX
Bkawwxe8KC9QxC1k45QZC1tHwp/GOreiiPl0mXSeND/4GBe4ZyI/gsbBzMpchgfgHoxu4vxKliUw
wzkTcV7Al3o5BCCH0Fqo579BLcj/CvLv+2yliJl04Po4sx37vHqokhq4tYMZR+/Lyv3M5bmcfTyf
NTjBdFkvm9NaupkH4Cmvn3Y8PTWTCQw9oVUvZ3y0wCs2HRi78k6BLK3TZ2pp0Lx9bAE9mAZU5CL4
NXGvnbZdGdZQFq777UyqqsYGSJOOBV4SDqs6HabkJqr+bUCIuWq6jijBBwyQpMkzjegKR1+8mrgl
P0AiiSJldYx2VgDbuUDt4R5I+sK0CB66zG1IIpmyuBXhL02Egs8K4VNHDtbrZVfo2o/64uWuROJT
OmzGFSV83BTScg4+NtCxXsvsq8XrfG5ccjluWgvw4e1dD4P+UEjpwzgg6/NsS/C92y3F1FCiO7cb
miZhFdzkylNbnm9sbhrCiuhMnMkuQ1RNRhhNhBnI56ZHtPryoM16dpbZCRJfLShFrxN/8VZZ2wcx
Pj9Ei4lhDXO2tQbrCsj3ZpgdXj9NiORwFRlXYY6mn0iMGtsQbyYLmBSUoeCPsiDQ1sKNgXphxm7G
0Jct5hUJuwGEGWgMDcbSjJ+g+c2oeTl4Yd4D/ylLEQnC5J/iLwx4YIQaPAsqzY+ojPVFoRCc8auu
XuWPnXKvfZyPAbKkfIRF/y2K6jTPwDuL+IuKa8YetKOB2sAwA42ZN11ot6mJg5PIlO2pTXj34j59
KbxoURNc+ZgL7Q01BH0XF6lC5rGvIIiJKtmTJuNoD9h55lP/RID1WicMOhKAVC+TTbtvftk811X0
v9yT5/0pxrcRo0IAA1DZxa1UwfqY/V45cfaTnX66zjWvpYUURIAXQYWmkSFxueHbp/pI2ffWT/2X
U3xMhraI0zbJKvXo45ccbmwweKIMIJaVcAT4dw1n1FtjrsY7+FpPw6s71tzd9pG7AxH+6JYM+ABX
IK8XaBUgK86mJ1bASUi6Qc1g2exxQOCZAOQFYr2pJPQAbAZV+1FLj6RqColCG5eFai3+H7RxMNaN
CFeCSMrOvU1CG3OAM2n/rn1Jsq6XYrO8kpR39pjyxoaQnHyL1q4JjnVEtKqmz6lmwJPOlzei2P9O
/fx5diUryWbs8w+Qo+9ld1uDjAdIXcFU2yc7VbMRogKn+GPm/xnN9F3WALUEv3mjyNx2Hwe/R+5I
hzvcFEIV8ObL9ukAHABKzG5becEeOl7jN6WuhIC/GrewTiLz8Two3wyx+zBRjEeZrBTMI6TW+SDj
r+kFyfzv32UgT4mV6rQUQGgQp/9MMSUbHF7jmn3I44Ldxh8mxEwawHE/p7dsIdSzveT8uqWLQB/0
OqzLPwhA/fMLhg0/vVWTBYl7IHKaYk1kgnWV3SS7OsskkLM4CuTVd8kz0C+Fr7DSpFwqJ8JqjtFh
jj6LE9w9mTvM8yDWTK7HS8/A3J5wfFxQVvUrbv9o/2YSLiZ90/SdUQVG2adr7BE918PUsB2ddtFO
7takM28paCGUzHUIxgJZ8KNQ3oncMbRuxkL1JgKXpbVlEB9uwGA5Zecy8fIIv5hmhbVKBg6jP9yJ
rsRUUO44OSsUqG1fnfKCSacuhVICA//XKRIbNjbWwKOQUTR/tj2LVz7puzidqNQEvAixBI+EfCC6
vvH5L/B+aPkM412WZ3U7tysO2vZkNxcogIP4vyyQ39akTds6GB3LwQ4mUm94h7d+ao4V3NX8ojhg
VXRlOY+7Mo2je8YFZJZLlUy2RjlW6MMKjaZqmMUXDWiDijLWjPHwDOwWt5tj3tmJqMnqao4gkM7n
AmXhjKoc96piZS7P9HFAjVz/UQwvfQN61Lu8WLTL4cz+h8u5ZuY0PrhB2G2v2u631D9s8SlCSYX2
X3jxuSMnsdatLphLlQX7SZtWEgVdNq6CA8h6FrMFMJGe4YtK5veFp6wEI53/uKqYVnVv6BQVgo4g
9oxgghUBPCH+Ctp8Af27/gle2SPkLHdm97igJJBZTQpFgXoLvXgCuu5sRivjvCrt0wPVdfUlEqHY
pFfegRgWE3Xt2LHGVEF0iEdR39Js9C/JlqlUfliIeNfScthtvPvjJUIn+CEmjKPMRuNsIWbN0lSw
pvNQeWulbsKJ+nhMQHoZPhyB7DrGd/MxNJXxFSqMWw5DlmP5mFo9Q4auUxN/IbU26CVh9KkFeq9X
JP36Ge8RwxoKT7npku3x70DOLUsMwaVwMQypZZ0JSiI5wKMpKoNrO9VJZYL3YubLpHJDIrgs3B2n
WAxNYTyH1AP24R1A8IEmmZclQlkoWQO2ZJX6OHMP3UVX/RUXmdFDN9Io2DuT0AbVT/ugnjtPHjQg
AZRpi6JJG4+fgJZ+4vY5M543zkIncwMjFNAhNy/l7FktefXH/4zYm4ngAbh/QNXqIymZGXuSVCUh
MAMgE24vrqcf7qoZvj9BrbaaO4Gn6CSG0AF7+gcJSKFbG7jHwVde2ofExwEFiRMJhgtxW37IZXeI
onOw4LgPDdXXjte9zv4vX24HiYmdnoYHwHhSpVdCEo58vyh7069NG6wEluz/WNTCPmiCc4C4jIuE
9qsLasfxOuw0YdRIu/+BZuGJb6q3IDr1q2RxakRC5OJLT2cV/us3GyKoPDcvgQhOejMkzIpI6nzv
NzC641BBOcXg69sVENdHwtv0kjgneXa83tM3tykHCStHvfRLQRVxBGG0WpFp7LRbfLHr8h0n8+i2
1QMy3eC8NrJqnLj42A4+qPsvBmEsGoOP3LEn6FpOl7bjAS3hFkC5qCbchSpr2JCWkAardTIpqGJt
bL0p8TnLR14tNw/9QQCz/czYI1al4k0jdiS/4Jxwv71HXfn3ZUq9Ok+zLxhMjFcpmc8uZGnUoKre
z0aJDHJlJbdyDeSCK6U013SijNWepEkiROB/TUzr7hdwQE37l1aqFZYfki2+vC8mO2/2CgurRP6Q
Kqt7K5GCi1mCAWG3TgU7Tnx5uI07CucYExp30kH16FUdblzfIFALFqgbJbwsY9qXD0Pdx2zWJkwr
C91v+5xfJK9b9Z2bjoUhW/9uNrhQe0dXWXSRAgBedAk24hUNXBEQMMg2IG4S4jREWEuVDT5BDHMz
C9OfCzjcMlWl8uEqWi4hNBrZv7PvCgbtHYwu/xIFowIwiavVU69/UPVCTCiYYZSORrIuGivCrws2
wfqRDi5/w2mSBiSQl4608/6D4StodXBVn9lRIrJ4V7CJf8k2OxSWt6pGEky/r3FnyxO+Xn2x1ffi
yJrr3vobm0JUWGWR46Z1QKyarI5cRTit9Kb9e1E2YLYnpm4jzjJD/glRNaSXXrHzSoE4CNC/T99j
+BfutYCInnI9G0u5/buMcoci9sjXk1fk9qEw+e+fRB+W1i9xHQHgRC5v8ScDiyz7YRQ5e+pN12fb
3VcdAM+tDWgSu0q2hUSnUrvXM0IgUD3dx6hAIHulq2qBN018uBFppBXhlZ+zrZ4XdPcmVwaRU+ng
y5dRdqvFE5R5zPun3Yn8SBPvuttTLkGz48PAecM/vz/4PyBhuhjlTt65SzyduJGpoeyD73JWd77f
k1xclvapZbMFSW+376eStiMhIcUK3R/DRMGLBgzgMzd6HXni6QGVK9dcsGtMajypMKWA116JCZ3u
qX1tQCi9l5HVS9h25qEMWMtpnLDI8ZR4hKgoGCwkiU09L94PO5MBZaE0kQSie4RZi7fEyyEfLFEY
XNlmAOC2zMZQC7CVyHl2ZpnhDThQ2l3vREBywwgNvR2d2wQ/iyIXD0XLubbk+OOUJ41Ttp4DZZyg
9PvoGxCDrTb5S9iPlEhOIfz4pSD/vXEtKI/qyOqXtbh1n/THxgrJ4pfvqcDFvO2oLdJcCjFO1Rgl
brjlDslT2e3HGfM6Q8asSWHzKswZYcRLFYuT4zEqe13fMnWAJ15z2uO1pUpp7g957tvy3xytUnM6
HTI/rLOWlKTbgrj35ctg8jg/skVcAlyyKozildPrTHrfujBr3PBkr1TBr6C6SPtB6mzO3wkGr2r7
VX/AEMBXa/wSvlQH9lqLMF5w8Nw+fXahyItZp5Tg4EXbWWfhYnEha4jW6lauGOkP6n9Rly2KsNWa
KuvWG2E3452lIEMEgHWXkYB418jntAXhPM0R3TjAP3LDgmv8aDehDl5R/lXMyBH/vFo6QybiOxdm
8HKhb6XBpbaz9blYJHF+tWGhjJrD95PzkyCMwjkYuspJgkMZA43mUDSgP1Vmz8I0PoBlnaK2/oP8
zwGCAcxFhSqWqGFPnG7WV17GdgXzsxb8SX+z0SaGFK2jtnfyccD+ecEbGMvgfQMQQoEu9c/GDgrL
JF2A5cGq1Frw+CxsM4YEevq7eVCOvIrG2lqRTy1V2oumN8o/z0yTHzPTvGZKVTdGhKRA2IL+TENA
QFzaxrFTDbqC40EBC750/NiT0/iE75FpSFzr9RDLhbbILdXoVgcXGhC1f3u3NChvIprMj9+OGbQV
MDY/NB1G1DP3PPk7JCGiqG2mjSemuv7cJxA4GQFwn8rj7SgjlAXQ3NKV95CAaU5M7iCjEWT+GSP/
GS3yUgpqybMVD0ehod8tSDCaaWWgAferwhQM0X4aOYVtI5cxz34psNJ1VanXloK5oI0pxG4X0Slv
i0IMDYm9y1UlOHN3tIUobalK/duqiOHO2X8curXVAw6l0etBERjjkNEgeLMWiF1TiRqvb/fNA88R
/MdfypJVtBCPorO26uN/CKbSEnJfd8+GqjMS5nzbc5aoOkuWQQP4r5qxr1bXmfnFnQsC+bR6KPCw
XySsiCqVyPeQpia+DjMe/Dd6wUzLhHsNiPFIGaMUBwuZbZNLNHOBhFuY9CDXxhBwMkSFI/Y2JHWI
QyubZu/XwhG0iWk1ndmzPd/q5aoNGt7SdCSiXw5EcJ7D14LqJua5nVar6EOGqPuya0LWCmPNK3Ss
9NYqbboED1P5iPtt0KDwuWFtD2CNWAi9EEo/XzEAAVEANWDL2Pk4s4Ho6pAkjwh4t+OsraWCm+aH
xYx/jfZiSRsXC8qDTTvR+sZZPnZXIE43ZW/TPhNbKHwkGwECSIgfZJu6YMKs6u34Au+ePWJXnBA9
7oSRCddeKah49J3X0AhfwUkPMLmCyPas1xZnsELmfZt9VHyPnEvu0RJronfcJbQwfB0FtZ8q1JLV
80T8u+gSGWfm7YrOXptQYFVQ30rtGKo7PoAPsw9mG11PeEtV2EFIMClk05ofC2bWvldTDp854tvH
VPCWNq7EtLqucqSO20fPEkLJm1qQYxIA+b1eis3M7eRwuoM+F+u3jSwZU14nmGE0Gr4AYmaDdRgG
TgKW56fbbqAecFJQsgli3Bk0QxSpYxNlnMT0ZXQbYx9KbRxORqtfEgfOEdicgR6+Y9P/1Ald1Stl
KR9/ynpJTQs+WSCojVf40gBjzsxcLiEIH7ttqI0F/vGsd/PLWEauwEz+Ax1t864tMROCb1sGhs5z
Kbfbwry3zunRFVbAQNv3fnOvDSklbBaxiYs6MgxVGvJ5zig37cbWjAN2JkdMaGelNhWcFXS+sBEA
KZ325v1hz9s0jDXCJsaEpG8fazjRZFnPo8ce350qIC4WMMEnaFZW/C92JWh0b906tRKZxG6T9aIH
XtgZ3dLUe+JJSy1qQCL9F0iUzFt7EXRTarj4bOyWrwGNMOwxW0bpTgVIWMI+5Tg4GNpfXJM0uyBk
+tRmKAXe1LBFUW9MVjojkpoVa7bFiISQCpeQBQsLnAMUoPPNE80VR/guI4vdbMBSXPZh9yatlkhK
CcHXM7JosUq1z2OuQQR1S51aI+rqKgSGa6/elBREOC/7JtcfRT8My0zrcGuEvovYb/ZujTEXeiPg
jhGjDYtHBZLFmZxfpYt2D7YczxDx0HFTyg/ZksdRCWLQYP+hUwbu1bRIYVuk26R+q7tOwYulWbb+
P9uPzF3FSjq1YJ0rQCMWE//D9PFoOnAX11JrTRXxcyq/dKXFI40DUiOpVWr8KgP2IaMdsPTqmJ2w
vbJBQtGuByYOrgkBGLNmpEeSeVItk/0IUU36XtXSsLF4yO2aXctQxLRszA5WGizn4F+/fY/t18vN
kbLbhiUj/9IYByWPP6VxqkTffgfijPtr2xVcOSzahUksVipxJ1fGh0Ec0/piTLgBwDQOZBHhcBu9
BFmj1MADsNg2SJWlNqg1eSYpQVQSKrSRcqctHeeF1j7kpxTOuZevKNbO5SQWifIp4fiAwlqm4IpL
rqgXpmEK3tP480iWMlmQzc+0CjBwvfegqaBouIJqorPnvS9MfHeb5Vj3xVq7FWaKl+AfIYufbEII
z+/3r2qwv8weQJorh9qmNkL3kvunTgrUymcKkxlZD+1BVVBj9d3pcm01Cg6yhBdXjkQYyTGzEoZ2
WcjYbY5MoJr+iiielpQiMJ1WN5GPDz0k0Fu3ytgF4jUU3AtfDbEKynmr6IdCpFGbSNXFL64E7FqI
46BtOHQIFcvuN1qKD74pSSpkGVUZtel1S24ZB0Rc4VkL8ogkLEY8HkQu3dd2UJFpy8gHwTiWqKO5
DxcXiul//YkKCk6GfhL1gMRfN6TxW/MDZXwLJfeB7ZMRBSvSrqInHYpAZXHyVOygbdMSXgMecQn8
OaD5xEJyxANn+zL2sKlx/HS16s9O2MpJ6w/e5OY2hVIih5fPoLJK1cIquIlpzGtJCHQehZBNk8V6
KMIbDylMYwnhlqG3eUn9FAlUmWRB5WAjMd0zC9ajwCb4z+I+nbi40pKc40VF9iZVWr/cGquGf2fE
XpeI/TueADUy3jbPN2Y8Tt7EjARRWBnWMwNOEQPKbQoGnnSNgiEmQNJg7WDOKUYQ9p3zWLS8BkmS
toB1AC/9Ie/RLKjN5uTni6vv9bqcCjAk1vQhmqgBqrHTrIBhp1ZRaMSzK4JO3puB2QMbx3oXx1t8
Y+R7CpNM0qSRwYbr4DIhJoG1ROuYw43C+frvHk3IRLoQvPKyJE8oaSBRJa4mK/B/N+dVZdbMlndi
yPdnaZtMfxREgU+/oZetznAAzvEuHtzhfbas+o8AHW459lVe6rPuinColBOF+QeAQVrtjLiyjhal
sc9qENn1nxgHQrqTvR3TXaZdmkblRLWtjkZv+IWFz2gJtbVHbsTG4ArW5rNROR+7LAtKorGfw+m1
/rWRXm/NqUqS8RUqZU36S07mmSxG9vqKIWUu6vEA1YL80WVGFOxPYie64b3YZFH8EkkEySayr6aN
VR2V7e7/aP+2R4Js3TaxFlT93WX9b99EYRRDrqCMR+4U/z5A8lg+5e2RgQpcbZzA7LCKt09Xeyws
1oXCLNXKuSEHLtsK0YiQI2Yx/avZtg17eZioLAyFAOhsPCqAVP3kntzyzWx/NwvurtC0i20nTHPC
X+zMaaA5OcAHs/ZpuQMi9VcJRoN3IL3tUzcTpuvByIo7XPCsw9uF/mW6HGBZMIXzCCO14HwzVAM3
IVSB2GHxQ9m3mmEKyQSjqi/Zyoni8XNu2gsU8960+VutSTqugzp7CJkAJp9Mlwx/BAoYskhjkBLE
6x6NFrMAmVG78I6kUceL7W9ahcB4qizvTjmZbudhxz1golJ9FomRTA7dOHdxvRXFsNCDzqyq3lu9
VisgKzvQjlYfudt5ZDgdMfQcL3ay/QBT/+pPGk1JCa3jnjToWEdGcvruZKGnZvcTSX3VNbOglEFK
WuHYUdXPcnwe819u+nZ439WCOJDbIUsY0FO/YwKyOpPfVlBKsj+qvs17vcHmSmA/4fq6Q4PZ9PwW
3iLKriRWl2Dm/owLeybPjgWxceUF0PStxAWctdUoLd7226vhY4fa7X0Cuj9StYziszi9Aqb+kcb3
88qXRcxZPbV8FJEuSeNF7U3znSWlaL7ght/Ble0vGF97xAFE430LnHDBPWXFDNJyr5d6TTdmUcLJ
5HFiTaWxJWIkpWtp4zlB5UvXfvPZraOgcBiSheSUiqxL1VPuGQ6uKKEM2UL9h9zlXsY1wIyu3jmx
lKKgnn+XmSj2C8DOMMs9rSeS1Zcmx5AYLGmHHdmbdfL8HHHJQhWlkYiOx8+lugAE8VGqltAUSw8E
kTvXwZ06hPkJMsAy9JQ7jP7eW8e/2RLxXe6WtAPrvE+7e4i/mVeNsL87E/ApB9VcC9MReaLpRGLH
kKDG1GEXZe7Ftlgr+gP9fPrxRFljisHPBLA/s8Tm2dgGBrbW9pHWRvVWTzxvcb1SBCk3nlnpc9GC
9WRChzc4/zkGytjpcQhYRjbSZ3aL4rc/OgD6+iqoexw64fRTNQ07njJ68SgY2GrfuamBgIhn6WBG
u/HmxJsV8Mu1KDWx0o2cKZo6Mm0ggJXtpgd/yB/+C//XbJR0v+FIYK2BA9IkR94EJrosbGsOb81M
N5cFPXwIk2o8rCbUW5TEIowruhK+gTN3JaG/dtt8Q54VAz7BATRDkXnFa5yvwzbz20Yx7/mT6+W+
y10jCELXLESrWOqfoI7CR86xKgeCYdll7aXHZQgihx28DgJYBfG8CBSJSDa4s1qJ4k0L91v+Od7K
CNcj//IVM5alp0nm3HPNSLX4AEhM1K3YPsA4wYP0GMByej/Rti+XN/ruprPS+OuP08IPRk0hK6SM
LPFOGT5LKHSSGeKy6R+Q9vUylnXMiLp9Q/1ZP/E61QUr4z4CTb6PPXgAbLNc2CcuDOXzvyIvY9S1
TTH5uG7ZnIHAFMYaS0/2aMF8pBRTI3LK0P925WVVDP6kdBB8G0FnAGb0Kys0zRiXK2fRjKTliuii
UtJKpOTs6a4TostFaHTCbl/g2tMANE7htIIj2HNuFQ77dZtXdTjCXC1tx61c854iV7elUh3ChY92
M8ohwkuIdGqwSuy2bZok87cXYp/4co0Om70tOAU8F16N3DITMOWxcagLL/Mtx+ES+sdDKuRBPf+P
OP7UkUgsTrbGvOY91aBqVn76hV34FtS1Nu65DrXLwcikv3GzC6qZxX6HAN3gQs4RI2pY4/IePch2
4nCvq/eK8ZagPIYG/WuI6GeD9uuGm7A0OvB2QSHwG22wsqGm1lkBBmfIoA0EH0QruNKNOcUd/LMb
PM5FP3AAxADBnSUWW+rAh2rAmw+xZfibfWxzDooh/6cdQACHSBGSF0b+kZrp7iLU/7QA98029p4x
WyX8mjoChRwmbeEpgEiiQPbIqEuvWPPKHCqSMfHqcj+xuHK1dMQfyJ0BiMWSl1gEdQJmJJw0ncPP
kZXgR7dw8dHbd3l8K+B2/Ffw0f+TNkW9DAIvUa/TgFVBN1AdX16i21HJduKrYebo1Kt4kz8Z/bks
S5zNtDJq2LfFrH79/VUxaqQweXyR2/zKm0fmVp4cfZN5HxnF8iZLHp3ucdbUdgRC8BgSrwrt6GNY
qwk2ZNyRSqyivBOXC6G1H/PU18YvKAa20ejMh6psmXliASp2ltSLBxjcVT+DdGd86r1YQ6IWTayH
0UIKwtMRy1bwLUna/YJfOs9YAvCpEvG2G0aAifnpcrLNSjyfPQ5ThgCKjq+XkH8AcNcuuFb1kxY5
Ktj+i83mVWuEe7/GIeF6Olb1cvpyI7/YPXBymjGgelfUXhMA/d87xb4rLSMUI9FXJx5uVE3ezm3U
WeTeVtqp/UxgomJz1owDeK0nBxgZXKertghLWhXx1mwGV+k5tHfkSheYX0bElBP7ebQTfpJUBAic
OiW6whX230AcSo7HGwLe083gfw+n8zRJGpYO5xETlkDam3SRtwag+6LDfp/aC2OYiFuZ9TLeItby
66TBBQniEqQwQjHNnSkQCTxtAz7LP1NT/aRxZNuoeQHFkBVHYgIWbrdZvNAQdAyQEad07aBI3Aho
o+wWIQOgGoHEAfWabIhJm6xTXfPASt1DN8zUxFRSwfJTbpuY8wpOdLcA1uzEFus0hC3I8GbARVNG
Z/aZtvdoGW64/mYceMcvT/S1ocEgWleyfS/gU9KLOUTnF6opUFeNcTM1t4PNPOlf5n73MbTto7dc
WizDBR5yBUvKU1qdH3LeVjDRI4n6LH4DqIJE3l6TA2gsnKbSliKXdpLeTyIxBw3vSJn3HAYW8LeW
u5e++J4mLm9FBzpaVWBHzqbyDzgodMaPicsn9AxV/QchBDyuIA4+kAfr5TLCF1H8gU9c63l3a3TK
QFaoN33HXrzAJBQqn+yEkLEtx9CHZeKVay23lxWLOfrBXKPx7T8IU0QWnh+Ry8ukMdN7yeyHJ9py
qg8yYdkSQVhu6U6YguPOo7hGHA3QroYZyx/qafswKx9dPIq+Rak0XUUM8+Puh1+YO32qDl8vmFqD
SZHOOEie4/ypdpCNA3Q2nkD6Fo9byYzUuK5Oef7pkcFV+/hpqjeNQxoao8zgg8Ht8/5TTWF/EmtI
71bYY1+0kMDqenh0CSxqSRbN7kRPT/Q0HFZqrce7UxN7D0j05iulvaOJ5zn60v4a/tWTe49zyQJZ
cG9HywS8Hm8n9LnXIec1zO/1hlBWokl7pDqaUu/4Hd4gbAj2RhEHqmegnnVEATqY8pls2l9VJwj/
ZTvkrZ+uuv+l9L93MfRnsyq2tYpz7wnJX9ZQGh2p2miVbkyKB0LqmJc8TGhJIdoYypVsp92u+csf
U+0SPHA0UzI/BvOdeoOjzJO62f/7CiDxR1a/qGuBG8uE7b40Tdrbr3JZ9DJ2nPEDhbPmwfb5kYGI
MkfRtmZToGRMc/lHmEZf/eCA7djQMvsoX/4UgNdCDGKroG1U2dABQY/kYdSnt+Whn1wGFsFLPKyE
OyfU0kcOi7pEgPRlX5QyoTBA1RRxbudVjqnzusnIvayEqugdEMnpc52UiKm0KaFaEXwyLQnOTO4O
7KmRQgB8EZapzD5nWdPmfOLfDtlrozxS+eVyg7+msF31FbsjLuln7o2Vdkb9VGy621ythB4/XaTB
7ksAhRjYvfxKRPBMMd1AOGicdPXcoh5ATpP33PkB6NIkz4818SQ7LgqZNvjExRqWSNKFtJ0EjWmE
h6SrgBnpPpVXw8LKzXteW+TO2GpxdFKbvOF/qr6g0x7GbMR6l1yd1MMOaS/qnol3UihwpEARmn9r
a9UNJ0ofrdzhXtEO9oD3lmtMAwlLVVQzcxBO2cA76jqrhdAIvq8ena5hIM2bwDuRvMv2uBGjH5lV
GUaXpyiRNt3hPFUHuEnJ+1rC1ErvlZ+Whi5LbGvzDBpXliKw3EIisGOPtob3niLnhfXy4iG7x1bb
nmWhZl0xKn+ROkALxh1Uk/8Oy+FXquLHXDqyM8Df3PraseSHcHm3b8C86OuymlQrd0DTL6NATzuz
0+SVPsGsVnv5KK4mjTpADl8mp/vhwZBnsVc4JytvP14T6Fnu1RVXWs3UpbckMhj8iE5f4GWJiW13
4nvPHu8D5D3hQBYI7GcbHS6ihymNTKfoa+6tfw2aoAZKjaCf2BU3gfHS3s5ZMU28FgPN+ufe3kpI
HWZEK9QPbnG4fZttcYXAce+MziuPIjKs2sU7x2vpKjfkHdV7FrF543zsJsJSUw8d9ZEqs1wCI4Yh
O0X6Aka7lfVVASMEyRhAT4I7jgJvP/30U1/gGBd3B2aXHlKUI7FVRBrnMe79W06AAoJpJFLLIPTR
kESgPcYpu0PMdcizWhQ0glFZzk7C+WFUWfXBQpLVipLAq2Zh+gexMZu7DhS6qmBRLPIhUp/EnNjB
2fELOJTr4ZQMia7LyMGRQsB87iJWHJUvIw3NBV+zd6KnOO0ju+N72UtqBwxYFthzDX89q8SOReij
12cwTllrpewDhRiRRwFSmJm52XXOQk8X8+4mcmWpMj7DaGHwas/5YwqY7z9xRNvHxX56NSB37RhC
Jrac26+6OfaYZEZFFLvTe3qxvL9j6l1SeFKMadT3VkPQKcow5DH6s34VaxOYI3VogNFO/l4Td3qK
WEP22xCtKXgJ+7BKVML/l/lX+qGGertVT9uLuX/V97XJ91xL31bgKdyqo3vvctTyC5bhQy/ZBHnv
uobTUZgm4Gb1L0wWqFVq486mN7ueTmPKN3MVQYt5LvPGVUSYgV97GvX+GDdFZFY1RSZwV5bM5B2G
tDIjoxvY2jLizaCwlxaYdOVijI9yG8etuIz7pxMzkNruy66xoNu4U8qAAcXAFZpY4SlaOAmxfuhc
z6fa3+bWqvE9NX7efwXzqNDHtAXBVtmbXwBxO+IKvF3qRc+edv5jN+97rNrcB+/OCLtgxe2XoghW
4RT+J94aevLZjrYhX2g067QE504c4lOMGsmsEWi8sz7ErS3YmraCSw0bQt2pctNL0GzviUlivjiy
fbJR3IjPLTIDFjqUYM1tWe2mSEADr55RxGZbi6AavzjrnQp/13jKrLFU1AcA7+IT684rATiY9oQE
/7n8ZOIYg+9TMRmVDIoND1C+ctJJfJQyMY/YUivq6qqq333D1sjtaLq7SNCXk40us7eH879KJA6i
2RA1VG74UesyC/eLDgIbi6lou2zfMc/aQDP2G3UI1ib7KuaBa9tibPCqSnQqMNFwJXtV73acv6aW
Mez9v9WDlTuMPps2EZu0uU4eFkYIuP78OFTCIwsPZ5eTT2FMDCSzvJZBcRYFRJYdKSAZqQjWIrym
omx4sHE1wcbgLM+ijriJBfqJ8gv8HG7wQ9/BP4YX39JCLroPWh9qSKHVc7Mx4wRCvpu7zMYRk+nw
q0SriralP2SIs3I/JryUvcb7rvegbJXcg8ruugbawuNBjM6efqV/GUDkCUwUGzNZLWFyNe67BtRH
zGXb0EglbXLK4i7Drh1aG1J7wqzDOdegTsmF15PmiCS+tiNPVj5kcHGVzqQmLA26NlmlV7pO4/od
VGDsQIHAT9h7nZHmjeAYplo3W/yHxz3hpNLEkh0clyHBvzvjEXXY2s4iavvf561x9oHJgVerzlLA
o5nf7FRnDAzs2fL0k2H6qD5ptPK7a/bzk5KvzAmb82cCsm+hq0V+QBCH0cYCCTsbjiyn6J1QhbSB
UUE8+7QeHdk5C9MyJomexS0U9SI7AwYNH0Qe65iPYYyLlweE402ZPBBpbTOThY0B0AY0uBLl6zjg
0Q4xCYbWLlwJ+93c+9pWY577yP8p8nOhKJnJxZNsUglwrXtVeqd8DKexXX0Opu7hJlIpX7S2S0J7
DoZymQ9mxZpSwWp4emsQbzSb/mtD2QQ5w+fKhfMrPEGnN5d7f4RDQ1At3wHqpSeDOWobvzdXACKd
tkv5J/IAP5nAh2wxk43KCJGsBhnUKr5IiYyWjCH3CqRQnnbhLd01mD/6rQaGx93UE7IUArTxaNxq
3ILPQ9C/uFdn6oQ1ohPSqFj0c3GLe8MdSCTCyZpARBxfahoky0mFYbuLEHCeZTqy6EzkniXvUrpL
7atcGgIOmWc+PzWZJh7w62POzkZWDuup9jaWZ6FiUkmqBgYSUkkjXjsGUFreOfuW/DiAt3wyThMv
2l/O/3eZqeSOgs1jU0zEhCsh1suTINO9SOu9uA3ok6NhwKTbXBoaKPYJbCMRKT7Bxndemh1KaW0a
tPwa5rCR7JeIo6D49Uof0tFWjrGXzD8SPy6Y/bk3mq1/C7U2xAMCnhaRk/+zxyZVmaOZu8CbWouV
1OtvbBlu2sAnxudp/QvsSiLJH94oKUwQHPS+XTsvGjK/vnSXPPVunyeGFpSuQAUAr/FH/DpTWt7A
HtN82OC03D/Wn0etGBq7N8pD8oUURYpxM/xPqODpzOfg0AksvZFszLnpcshbOIZWY6gEcasRiO2z
aPUfKlOv8XV3UVlMnvZkob2L2ut38eoKekrxnBuDuKB/67spfR5gpgizRRNttqA/V29cwsuLQnnv
UOj+dchBUKYTLMLi1M0/Z7UWhmNXWH1lEBbrGrgNsbWmfVaJl5L2bOF7W9tjaxKDna2EMseGBEBM
0sSYuzWWZZO/RBpR063pI5iimgS2C+yCzV7B2X5EnSdxsFtxE1C/mkpcnKpk2knDO3QGfWtWRKVI
M4p/q4Q3UfIm28nLwbPKKiFF9epse6emZP/UOQvluDd37b15rnizsREx9QQoD4MsAKoH0rV5wMIN
5DzXm+iSYn3sGOeaJFBf3ZHwfX38/P0XCwzybgR/uh0A/bDxYRfWV5YQkB55sAMVBRGYAMZVp0s2
7F4xCB5O02Vz7HiG7Aux2LhEg3953vKbFW7FcchtXFdu5pBjCcuFTLHAEcVxc87SwyQM3N5FTpcN
ONgPJyonvENrAZqvzr1FeuIOdco0ie29B0vdbBA+qLr+mfHPn73oAfFls7BP+trNaCp9mcVqx0yK
jSOiO9Aem0wxS8PyjdTnlbj3svbzEj7I3e05Ptjyv2LIetBoAQZ6EpQgP+z87pujQKmRrf0h/emh
t0GO1kO8/1Pvh0X9bVHCgr26iZgPCPOXIp5oT/BAXLe5ytzZqb6PwvS1IYv85lNqO9V8Tgj77vWA
nxgwhFR3lPJMqotjeMBjsJyjOGVz5ER6IcP0NMOwBCH5TmsTUQ/TMcnV7yRghzhMSkxbFDcqIZAD
shBVcPPkw5TddRTG1ym8B0FAQ3nxJqKjBEfb2d0L+bSKzZ/lq+6zsg5B4n3+GgQbuqYhfPX4Dxao
QKiQjTu5jxW4suCJ5IA38GCtT0ui0kNFfcGN9844uEPZi+p/mkoZGBCO/63qNJRXdQcfOZ+QRJXk
SmregHqaOru5FIbd/uByHEG59UrtkObb5yLvzP6Tnp0IbbmCtVMYBfMeuabd0/xAL3q/qIX/PFAO
7Q/k3Jo3DuRa+K2vGxpyrUo2CvnD9DU4rM2o8Sj4ZVXCl5RSfpLEPTw4IKZlWmxabm5vv+6LNXOQ
BCmZnStAUwt1K+Trqz1H1hsjR+3nonk+usCieFQzQrx1RX8pRD27bPZWtZBze+HYps5iNpEIDMRN
lrIQ/gCtW3CtrnBHwT3KoaHIHy2M3EUGgnypAgPgATEILiFiOZM7dsUTKtYjlMBOf71aCBf3QOPR
PRGUeJll9HowLnmCsPshg5kXjYobRkb6xCAV0L7g8WpZ6yKzR6eUSqA425kLBfV7quF1RstXKXKF
74KaOwUNoHL6V04Hs1UJCkkdvicyFYIRyL3IqYLz1X+phGe2vI5tyNyn7tr6V+J3ADU/5WQmVaZr
JI6ti7SlgDzJhKxromKSYT6ZoOrk8JXy4pt/mCntW+MQBzrZ5ELzJeqZuRdSwvf92I3hu2GHnRAB
Ofl5VgXLNsEK+QioEiRMcyPPhcnpuH+KQBk39LIdeAp/a51vegXo0uasJq/F04vAm70BQx71XH+M
DfgL84REScNGRTWglOAgY9T03qYiMkG/XjDwmOxKVM5cS267tdq2KIhuv4gCmGdvFQvbFAse7JZU
gD4w/78HXRJJEAGLaZeVp+bq5jw2c01eROvih1z3c/yyybW4kHyT9M3Lz087eHsZsFwOia23lzA6
S0Ut9BHf/InRPgZlV8utqYMkzbeem2Wj9dLaGrC8dJDcuWrqi+1mXnWO4GLfv1nL9J+XfRXgXiwZ
DajUCqUwN9v3qLGF19S6vrxiAEbIDzu/VkloCC6MFJCft48D3SjgjsdhLVsU/Sv9lkkf2wvxZbLa
swUqk5LNqfyEt3WWS2WNg/G5h3oO9+e79FpODSFVsqEj0FmxJwGK/juee+j1NW2/Cvhw+asg5/Rt
hMI106FpBMMQae5fGNkcZuU/cQdOiFkEYCs4Ur+a0KeVPAZU4WQM358o6JXHPpdJDIfhASxlmxH6
5iDiQ9yYzLGoQ7rUvDFkH/rBkLvE69mEREAc+k1jtrd9S3lj7lxd1vUGYB9mehRDxomOb56DL87b
LJ/zxxXpk6+81j9AkvyrPA4ZZS2OaJBzd92QY0QwG+ZPPxFikIOVHPqc+DpyS+t3EM1TtbB9m1Ds
T68xNspLSB4AOLEekXotw67TszUSrAXzMmKXgZwf8FTIEyqxUVbsyiSGe28e6eDqc5SYAqmCEein
Vew127fCRcEMCChRnuK/8bS2m/RdkBnxuf6z/k2OU0FrYWMGOPPOh1TzKwRAK4c/IzLLzawxQ14i
0HV6gQzA6zMn1TCbkKBWVfj3vASA/zcULoKjhumAesIbzbRLmEB1ZbUHIQk2zR38ZqhVVF1bIZ8w
cM6K3//EwkzAJMboGtPvRa3eeUNEW86fFzzT5k4B1jD2hSYmqhiAi14Xn7ZkjThCIOA9V3pSGz7V
Fl0ycTNdwiQMKRjPs6OV9LYyu17pcfIS/gollFRRFlghCutavGWUdn/clcCOLFW90nTx2XupnBNj
53XdGzjkgKljyFIonpWJM3BlCFwbp7qyjQcRrxwUOsuAHaWangBg1bmg6LPHWLvv+DWzCfyg/XVH
3wD1GvcguhOLD4c++4VL3hCVCPqLvcRJQteO9qUyU2pAELjbagaFLyVi32aWARePgc7WDYBA2kX6
mqoaq9v4RNDPcJczxLla37Vq8ifIHfiQ9Px3NKNkMgAALRtUKhdj/mahILloWFmVF37ws/kr+qT+
h0ZXlOEOKLfMeSe/VNA/rmxY/gcJ4dYTmxy5K3HIVn1trKgIJgSN4g//D0gCUTsyoLfG/U808yR4
pAQu+/MkiCbYi+/7oE8D4IGkzVAADJp4YqcgsuwJg1W03aE5xWWCwDSgsnMBeSrcI4Hpg7Rk2tnj
dXI78rlhFJwhUynpEFilcuMjMi8N/imIVa7TnL0dAFyoW+YoXuN94CV2FkwsdmQo5A8K2+xHewGN
27Q9koSJXxW4OdbceLgPuMD0LOQS18DzRmyvlXf1HSEGFh5occ9f3xngpc43JuOf45dr6NPmus40
6O/jbEwYy097o+JnACtQhkOq4xGKg/CHuQPmtirh35hDY6eOI8QbffQV+iOz19KniAR7DZTWPExk
MSBApoQVc+rj9Qe7SyYa2/61kWB2SVC9kkTzh1Ajj9qHq84HHCJCCzebJ9S5tt5te4PjTWlQSUQs
gv/s11NNdicpGjXc5ls0poofa4FG/FkFRmCEZdcq7wrZ0uTK9O0heljtvhatspWRR9lOIDQ1E+xM
zmwnvOyXVBKTNHXHM95CoftTH/dy6ZiED6/2sl93gwj6qibhbtUD982UODKAKvBK5i0UHGPtSL6v
45PGHmULX49cP+EOUre2kHC9nTaxR8vIdA+J6uJbxktnGe3ZLbQZT/e6/XoGyxiATU1gW3wcbPEO
XFkfAr9eoEinGkUb99fChwhqhB9qB5Vc2zzal6PDyoxRcwTRJ7Fb6GoS1vz/SiUtorEf6gRPfHEv
DdCwMACQMVzG4ZuPHvmrzR/wn98O1OoWmHYGZnHjQHuFiQYwombQs1pP4u0zoh/Xh6O3BhmZCwM8
GPccJ1CoHkB76fZBrUBvtFA1B96/hEXUNFudcW8y/Cli0Pi1f26UtriBG9gK6qOvlBDyCsleqaqV
gnwbyoIEubMM2CXtkPEocoNfSO4SomrevFHSZN4Xa9UT7PcoDczCAB3KV9ChzXlTIFEA1mmxfUcn
7M5cb1ququansedccxD0r/oX3YCONq392+dukR7THpYiUNIaTuQ0JuADNGHAHtRcfMD8BmrUCUao
pN1uIkED1KCXe5/SN5mhEhHduvh+DDggse9gTRp5gWgtTC9xOqpU4EPCiOhE5RtLC47j+0rz6gSI
qZ4wzIwxAOhrJBnfeEIChtCn98wQmBXRpRLb7CvbpNBVWbliF/rpEgQaOU3zsM6OHANPCCfByEmi
iAqvAyIeAYhyn0XjbwoHgINZVKXKu5wcsqxPK3lvgc906jCufiGH2zL1HO9G6y0KYQ8k5t6GI6E2
UAGc8Rs/sq7Xb77Oo50IUBtYqnvvTXlKXM1+o+kpXKyhnFsDg7WvaRik9IvJSEeK4C+MQqvcREUl
H/mbNhdMdsoPi0+6j9B3pbGz59nyiQkZQ/FqkhBcsciNFiwNUSKdEaAMWU1OppEFtW7F+zGplSVO
N72zT03EB70DlyKQpNvNLuTb4o+qr+SME1PnQvOT26yyTrSPEhpaQG9FtI+bjlq7MrDz2C5AuMWw
rMaAOHjMksnnB4R06VHaFNsZfS0HTvGJ7YHcW8LCstLlA1VNQdRMmvwA/8CT7o9ApVQGC2p9G8Nd
yp/CP60hUkoFli4+a3FO4pTb1Xm8wFrE6J60mbGVLYIsRrc+MlBBxY0lkW/vtxCLO0ukF2qZnwfz
sRW59+ftmRS/taY3dn8Azz9lACEd61c1abiAPzP12zBixZ3yIrlbSe0pgFX7rX3KLYuCewIsHISn
ZErdiQjXWQVXJXgm3Hmay/jAEYBiidsZ7OeRB19kQwM9Rb1gqKbiR1ZBBIFy6bklMVqXEmgQjD3K
O3OLMYztlEZ4iVYkbUjQ9qr2xjHylnmtwoqhPJ44hwRf4/jGCnwF8ThcXPJaSKWXQesp4QTsjwb3
xDSd7ItQzynZOIToaA7LzYa0n61nU2xAg4BXcEylgAUV7ss5NQUX707LY4fLzKMBFLtqn7frmd/5
Tg/u5XudHk9G3g9CbNwo16YpVWaCOSQSkRbbJrlY4X6BeEGr5c0mhgzX96smLJCxVfHxKFwJVz7e
2kRHaVTVgKdxDjvTZW1C7b10trjXEukJDHQgfniGxu9/25re08orEzQe8QAvUry9DNBk+hR4cX+7
c06tNhlXT02WapRbu0xDmsjkqATY3zhll7aTt8r+Zx1IqowwolLLDKu/xE32YLuqf2voyPfg/0xW
2VHpJh0sJPgjw9QW1haHkK1mkp/Ib+JgnXmj2KIQcZPL2qWEsBiwjgSYDQwqLApt8VYrDlnHL9vE
QgHlQNbm2zEJwaVy7/pT68qpWO9He74gXMgwA4fSj8MqXTybcSiTbCDfyPtaHxYQiZ5VwznHwsAJ
Xwf+eAnUA2dtUuMRYQbf9CM0PCPI/zgV3YGnymOfmx10XfYdBBN5SVmFaQShTM8HdOdE5vLRU35S
+auNCZDjsajNQXWEdwcfpHfHQW34yJHseoAfI2GMq+sC7spUYiYlc8MufXrGw7RHA5tQDeuXOT1b
NQQIJ1X07QsrVYHs3bRU5nvp257tpeo9I7nxXC0bMG4ykqRjR9uOZxud96FPQ1T71rHTKwkWWAvo
YW1c1jsaOgMJY1M1AAq8ImOdLIAq9x1xEE4OOqgdOVyFFwH0N7gNgHAi8/QZ+UhWJQB9tc0SsALi
2HWylq3mnFPB0Qy+sWEss6RKLdf+9aKD+rIm21w9CWtuK8D4XIZH3ORbsUSem/PBeBUTz8XbRPT/
tf3Iv2Je+xnb7ym6vmmH2xpD5DNbOECfCO9atr5yb4lUBnC3BipTldAH2IQzpXN8MJVHIzQ/m0UC
4oBzXRNV28I5z8kSsdib40tvViwqKAyQnIj9aH1r/9hrgISaiYK2I7Y8jHYc6mAWHKmus77ZbyoH
GAxnzZhcTrupKJA+151pXJrI4wB4b6sTyVqC0sSr52yPtBVnTV6ZzvJhspBjUd87n9YnsuMryYLj
NxBvIsy3dlcdtKFy76ogVZIBlKg7ptY2SORlWP+pTLP16W+7lX63JNquTm1XeKzfB60N4CAST3Vp
+DiwFmlwgRduanc596jvj1t3JXqMNJi3e86Yt+XgnuOJNRIWkpl63+mNGrdKvAtyAIsmRUsBCR3T
0p8EcLwGXq/FSt10ajHp4fm4SboFPwbhZoxczPs8AjBLzAHrYu5A/dxL6sKAP3dPUbRGRk6mbkaB
ma7sDUB+hRWIcgaL0lET1cRu70TUz+8DhJcjoAlLcqX3BlKjmzIS8OcNfzCaYswKd0dOuyLpUxIg
dDmxSoAXJre2eSKAWuud3vtm3iw3Z+bk02ILpv8XHpEmM/860JFrNAXBXpahgoPaKKMYTlJkBfFC
qOYqZark/vOP7Gf2Dx8b6HgSgcZ7IR3sN34UDvZ3wLPXuecf5c1qq7JPTL0W/Poht0Li0/RXGqYM
6t5hRuaWH/JI6HBEidvHpSaU2HwMa9c1eTOhAlIPysQvrnwZtlOlF9b4Iac0ZU6lYTWHTGhkUfh0
/OcA0lEEsNrqZHKNhJKEn/CPsYdVzvD30DAMfvTce+fm0mYxrGgFJKgfVbB5piIqQF7EOOYycLGY
Ui+50XWklLUaoyMGCATrNOuJfQYF+T/veEwrgHCE3tlFASbPwtuSdWH0ozISU64maQK3NpDS9Qaj
01jAEPdYimjqbNj+BUmZQqovGSBx7UifEgFq8iSJ/Eax5AZQwcEUvbjj2CwjB0Yf2v/kWzWT9y91
3XUiecVWY4NMp+TRPY2h+p7cNdez2S28YgtZPb67E0houJ8999XicqnesxULNjrAg/ux2LyvAaaP
IVyM0rXRgKmC2YoF0caG4+TW66cZq4dPeCYxp22M9KSZy9wXqsvARHyV5fwmVji8xsaeXQo71ioc
SvJ2yU2ctCaloiKho5tzR8EcxUh7R+fWfAGmLEKi8uzJ1sprWR2AIWkO7PHaWQJIr//WAo4LdKZT
GfVk/0mzlmmvtJMgk6NrVWrPy99y6zs8XysZV07XZNtrI0VokVG8ZO5sDBIR/doJLHC09Bfdmay4
fWhfQUozksL/iHrpkln4R6Vdsk5Q4TwOUXPzdvii3arMrWYxIw4mkS4FSh8pQSdgp8DSbbhgY0GK
ytj+Yk8gHbLH5shJqjnyx/YpvmrLy8zpyXepy5zSGWSPBhYj4SjDSjhafgWjHOuoxCriRLwIsMFO
w6XdvUgQleOPfKZ2SaCsrO40eSrDoCwLJVTUARVpKKSuElcJbZ2eXCAqKM53fWfk0k9OCMViVrFq
HlAtd4jPp96Jl+9M1tAKqWvPvvkxCAxejq6monY3N0n3Nle6u+zeH1DGSWAFhqMlD/aLRGAFoHnB
og0buOlBIzWTtGXCsoF8YpP7/RO87MO0D0Xk3anP2E1cWmA8g6EJeq4hf5ozQtYkZf5dQtV73pp4
hywMveBLxYZx/7z+Wg8SjNf3uXM7lvgbo70VJZ92DKdEbybKeF0iLZXbdnOCyllCc3CQBfrD66kU
JF9+IhHlHsRF3xGniJ0XyP5R2LByg+RDVkHReM+EF4NoHr4cOtZz2GUnHyYgc0EJ8l9hi6Ew7k4I
KK2v+nGfaJ1i+TmwZTX5hoV3PcgKBtgiw+uo4+6E064aEIO9tfmYETRjONxj7lCGqaN/3VqNEeQT
Pa54nu9E6bcIkiMwKupCCP/hXd5akb/Vo0CE1nInUjJpTW1+sTfDm06or5Dzt6LpDALmUsDyB6Fx
quiTxiwb0FYSqB0uQqFeyFK/VOWuudMcQzXQXgygRxITGduF/k8Zk/5Qc1GRuT++siv2TS5kNvyn
s+7NNxnVJXkrILaS63ROS1g9he0Qcsv2Q0ncz7kPS3llUoLuYEY0gleNYPdMoLGdxDZIp8trgLxQ
OljOgLczB0xQtytqXYE6dKpUMhWF+92mLVYAdvPUzi4LvJ7Ds3DNrV/RMhvjGPDGpo8n4P9DahfQ
T/0yC1C+/+KY4ul6BA8T5AVW1Zd9DmsCbzxjNVhvCDxtGK2PmsuEyyQNN8nCt7IrrHz2LCq2pPEu
q7z5C/0jADCekBbnQTASTe1l9evOGu4CXrr6PQVAuDJSsp149qVZjxsZWOa1lTDOTAfzHte//68l
oArA802aXXOZ4wTWEgLQYfKG769Vu7N6Me2vgVcgbcHrHixq+EXZticOxiUvsKS3dE0fg/uo4j7h
5YR5bMU8y2Xwvty8kLdYKoq94nXlt0ejSsDjefJosFS06mwDyKqr+4LjAAnH/yAxREKDvSEHuMge
wW9Sj6+aCNqtwqT5Y1h88xilEp44hjAML5CxuTZa51czDDqsBah48mDXqT7kUdxrT5geXpt8ANIx
km5XVzc7FR+8G+CD+mYcunBIUTEGqRg9ar8I/cei/aHAq6KCeeyAdd7ld+2PkFHzdMuO+LviVjF+
zrwaz4lScImDeKfhF0F7UtdBwWTg6GxNswKbNSRvPqs02Vb74L3iu6gMGuRI/sEU+yowyzf2FKEl
0HEo8cKSu7m8i6IT/GnKQ5mFdOOgRWWAv33EVRASp88btnfS+KknILWl/b45QOQ3IPsGtzD17GA+
v8YYvANAikHUgb56Lt1yLMv/yY3z7fu7yVh9NQL/SDW8KU3nVj/KIxsbNwmscV3Q4N+aWNurl8/r
gKcOO9TDfkhSVN0sQ9zQxLDCwt5djPoq7Db9Zh5Y57qKZJyTDOyYoCUxpnrMQyxW2W17Gh8M5rIW
s1b2E3LYaOGclrzRvHumyQL5fs/4G0qcXIjSYDi7Iw7fPfoYvlWFaDeJBn3VgOKeN6DXrhWKmiGO
C/6/k2RCudOUrdReVDo9Z2yHVqVTojt1aAPh9ASNdXl5U0bLGb/AK4yko0XARxI2Ze5YHzu1yDNs
dG23wH0oZbpAD31swMZa8gy+n7vQ56MVfBslgyJ1G+D2/Yi/qhSJ64DAfnwYrRBlg+euaXjxqonX
CtX92HEXMMmdasHK6uYC0WzU3tNd5UzX93S13P6tVQK12eNLv7wP8Dc6abT9bu0F1gU/CzfPe+x8
smOMcdGneRdnCDw8LMue+bDSw88X/Oag/6h8gpnEVxubTksuI/EwmYBjFgaDuyDIDBtOQxDLkW+l
0V0F8pO6bM9lJ8IXTgHvGUphItOJW+b/GdUKT+eRknHfqzAOt2syfbGzpqC8nQ4wQ7rr4F+qFwmx
j2Q2RS2bceLW1+UdrNBI9IlsaJZEQR81vPEVrcKM6MqXxilCWMjW8jdiZh5XitbGR35heyA3e2qi
HEMvL5DySFSnVw8gkaD0+feMHtqC4RZKT2Y0J6zei0+SHiN15UWVVcfiGJGmJ33iYI6Pwmvi52RY
vJAOgwus81KNSEH52WjRn0SJOlM0YsM9ea+vEd7fAzaPa243GWJZrTmhkcI2qBT6lH+veiDwq0WP
XZLjPhuRmnOrWo7EpglF1sBwaGge1oqXwTGfiecQ1O7+peXuqcwnAc+N7GwG1hoVGb4Yw9iTVuNz
ptwgMDuMkcne9kHR7YmI/tW2izJdQtEmhvhdDtLuIsOozw+FbYiQXlBUHbLpAmrJoKDd2r7sOkII
+eIBpL7B3uFlseipABM9jtDMCA15Zjy/76hSOtCTxzGxcx5n6FlFExXVN7FVOCGcHPbaB1GnWPLV
wyHhcAv9mVnTycHNNaK4LD6En5XB/LgJmYS3VIbQSwAS493jh5JO1ZaTdoRtj8QKmzVKlCTpPpsa
VPRpI7YtJ9RP1G8HJkyYdavnwmSOczISRtm3QSduh1Cx74XRReK2j/er0f5erBHFa24RVwv1/O7J
bmAppWXaZa+GgabkF7eN6IP6RaGHM3NaGDNDJwnygk1Sce0vh/gkhGdCBqNF/m6a7D5jD7nock/D
6pacwioMuE0GoPKl0QSKhVvUB2cifz7ff4xX0nvPI1+vjVhgGxf7zbbSsW5ws7ex7vjJ5p1DDkS2
U9/aVja8jK05WqCK9UdLvOdBRy7HnQ+ZI90WgHNxutBnGQ4DCaYQpG5Fe+F7q5ufGgObbcQ7ack9
vTV0ikCocCbkQQEEEOsX+AoNeE6VezUP/E5U+wEvtU8oprHiFBjCjyX4+F46iA73tT65DoO+yS4m
js0i56HW2LKcm5nBlYfSZQAdXOwDuVnOW8X6TeEUy3qM9TgSPdMadIrX1tUtXKxvyoS3yyxRF6CS
TlFXGJlZbpTkRldr38HOfgLNwppmopHmAiUAJDq0D0UlnN2ZD9HVCQProCWeaLY3Bdu7jW5XPxNc
A5C/JyCxSevEv1gI9lvyqQnv0vrH03sHJcPQtXUk0pNJnpsOnX97/rWYoElw4PrprVAIU1TV8HyJ
Mxeto6gSXS30iTzZ+lkisqf+mRs5EuC4jsCzkELNrX0nQOQB9P5uVk1+gu3y4ML4uoWmYgyXGe/Z
9RjtVWRQ5S4cypsmNv8/KLAazaP1sELp12SOx8y+P8bX48Qr4PriPNFV6BeEO8B+uOctfQ8G+iUa
wg9g2jXccdfnJEQyXeE72gpdwj73pCv39PtE5bHsO3WbjAa667uC1bih9v8fgyOF/xQ4GMdLRup/
Ud3+uzuWmY0+b2SzF+srZrNC2pqHW4knQSSuqeMUAsbLFtITkY2q6wD15gTuuSpHyQgrVnxzJgn8
JSu6BiNSzdEO7vabGE1eMDhloIpiyIyOsx+2P0whI63zR+g8yyIcZfi2v9G3PjTkhJRSF811iWRX
TrvgwCvg8FYfVTwkc1BfE1tEsIQ7r51Hrttb+NkzD/AIt2KeXFsXX8JMB76XB0MyLMlVe36s1/hq
x9WzJYXeJ2Ggb2+D1bG17mxi8BWDLp2Ffd/unRserC8+/TtE9hnmj/OUaFrTd6E787sau3rKenTL
OyosI9uMdk/XnR9Du1IowOd3LngzVKESI/T/9jUoLWG+9ck/z2F8+kddV6f8FFpIajQk1YjAPPi+
9eM1Pdavp0ycmVxfZMa7bqYxdf/A0PUeRN4uI2OvapGhN+iwG+/6FeEfhcwTmSdF9n4M00qogiMT
PPgOYJ1Xl0TxjyhIqjti8ZhgpWj+vsgAsd77QafvBvzHQo5DuWL+m8rYoOwb6PGtd3Vefao+Sj2z
5XapBGwjPX7W9478+kdQaAz92hlpglexsSe4pd2mEG0h6ws5d5agQy+iLBkMpnhXoPi58la+FvyR
g1ugafm9dtCdbJcty03Ed2rGn1wC3Q0DtBLO+e9Hkv43MyRGouTl/eYgs2zUWhmiNfM3LtlPSAC1
Bty07WPr1tVPnvAY4mBsfzgpP/98mMrxcc84RM+T5Ep2n1NudjYOPEj0dceUglH/OZ83aNAyFzv8
T9pFtF3nmBG2VK6GpotsG8MfdjFNYCV3EoHQmlSWdz18/Jw9LRYwzkOBFPKq4B6dLKvFMkM9e4ma
3jToHStdoh41e8ifKNZ8uXeoeD8j0GU7dAy2nymlhIm4GqCalRlpAuFPH2rPcA9D7wLw86VVkrAM
NMTVhNG0GD3V/0Tf2NcpEc8IdmtuZAwFK/NxcpZaln9iVy0hTaGtmvkrtJeZt5iQcV+EKqKOXTWk
RTWyguKtdIb+8Mr/t3agZj+V1xt5C4txIoqpAt1rheMuztwXbxfBOApaCmQX7LgFrcpE6D86g9Ju
b9mAFkGyHYgXpNAHaRp3dGQ8jAPGiGM23iPH1HlSwBKwTzeP5GL5LVQ+Q+UUXBB20DsJrSRwF28R
Iyu1hO0oer+TJy9dJ/EJC0VYr2rkHUC7VY5bwgG3k9bkmTJ7QP7odMP3ZHXHUoZnsmvEy5E5SKv4
rssoAra0E0DW4SqQsFUv4/6zE3/MjJ30uDHDeZaXsefQmMUQlw3h555d5wPKFYfyW6MEMrffuIDS
W4r4gi02vWrH7qAgCwT7y49TWOrwPhqDiqqmv4/OeDoNdF4YupUq7pFOPy78R2I6yhyudthy/JG6
MTBRwo5tFbfdL0IwytIsOCxlg0tBOpxIWYHXVADik/OpNgnuxABJJpqZV/dqdvIdlSZfowOWdJ+Z
e7QS+7y7FEnd6giBw7O6OtugtxbKrMD5JRWAtCCph3QeqtA9S9OnDce8WnN0z6NsQvqOfrrX6/IF
Y8wC24EaDmGW3bTHHpk79qQXgteSLMLUd3BXP6//kIlmvgDBYqWtbGUmdZYCExhrG1LbNbXJsFsQ
gVCmc8UMUvvSR80g4EtutyMRz+4doCHwyLGPEPvIUqmS9MJfN+wvzqoB9meuytWzFfFuz0KmHMoe
IMoPhrTaKDPswDiDTsc9HaPAz8YcfWoFB0NBRdPMakasqtnLs2wOb1US/2cZi0w3+1RsJk3HNF4v
Rj77eeNYjkD+1VVU4oVyvhViREVtE8sH7gBZQbzgVKX4lTW4YGx+2N7nt9sYdW/Q0cSx6dbZ7UdR
qvh78puTG6MwLm19m1LxfGUVd6nuZKp4S+OINUeoipGyQDROl3lO0fZavLB+HMJgaFk3s340SuaS
pYIJIN+5A/EqYjeAQZ3K54bC+9/g6AxMgvIGaNjnf52+rU5FM+jU0igoTa7drFrnk9VGkA4Q+Vpe
//1XEqcti+NN9BrO5Q9P78KIA1rDh/bcDdD/gL6pb77aXR7XyGAWTXlfikpzN1XR7h8+6pp988TA
ajCmuGXTOcYZlw+I6coEw8bjbySyM4o2ehS58mJPThYQCh1JYoxWhBsmc4Woo+0DGZgNgUGGLieU
UjvB066+T0V1SucRAk4v83xR2hwarhc0LEr1IAsT9+B19fbJOZ/HSaNXilp0GZjW5xYx6shzREpm
GA4Xfwta1DUUaQMyxXk9bwp7ZzgdzS/wdjxlI9w+kX2eS9qSIPmJOicibohHONrTJiGcpsgwOI6i
8thiYbWV2LUSTkMeK3hQS+B/k7NR4yp5131TmN77hYMsi5nmg+q16Yp7qckyMZIxnoq+OJ0Fqg8D
Fx6GWthOK/PbmnrufVBX4wuZII13DXnNG1PyuN021f3W7jL4N36YpglgMh4qSADP1TLbBAOMxo+1
OpnyeuDD4zT2YhDCBuhkQWY3vjYwynKTAyc3inv+dpW3Q08E3TCb0mu+1g3ZHkw38iS37AxCux2R
MPTsrEaKj6qw3cIfrOFFK0zZnhrgty/Uluw3GuX04P+44NoB5pcQamGfPa6/VoDggtGGf1UdfePz
oQ80Khs5kR4NOEfL59HkfLQkp0M1wVNkdnSzaZCjLcTioSkJHrJTfa9lLsw4wuLR+hDuGpHx6o5N
HqxUwh1KJtEmCyNXYe7xR/66CKV8qE4N9TKsRfv9l1U4CUem1ditAZqlcgVHKRPpKqmuLTRcRd+r
Zob7lstCxVZzuwX3gx0ZgK3fA2e6jV6pbll38jMW225rz1gIOYT59kYvqaqOBUjbqEIe93iCpUxM
BKqvXESuP7UeWBl/ddWjW5Td1zO708c1e8Ly8O8KRHVIgfXkpRyxEL4U86hobNLHzqZLWyTispzL
DOxltrccUBKOQSsjvStC8TffOTDP6/2puS9oU5eEBNNczyiE6umicHMiImMgIwEQlQM04kce3iXt
GblRXH0zW1E7mWjnIzw67SNhT5tvd6b41DksPZXIhfoS9bRsdvsF96ksZyyDzEnBxqDYRzWYaSz1
6YMeBEL7lKKjX53Kxqdb3roxVr7+Sh9OxiqoUJ3AqRJyS7yoT6k+pwOCXeGqKes+jG+MpZ9BdJ/o
rvCYY24ktpNkDhfHm+BqNjJxMzcwUgYq3Blp/hrKbN3kZIsQ1e1EacXwQbyc1jqwdXNRYypULOOz
a/mZn/eMwAnayqMxq0ZpDM3TeI/fmahivm+Z0lATDSEuUutxticCo1C7vAAjCmnLPxbRJNBAQhyc
8ViqFLoYfZtGl4rNw01szApDRXVZsNVNtfTG4KnvAg1tU2cX6AhypWcrsiBXigkBhopbOGXJDDiV
/G9C0CLYp1ooU6s8tb9f3hI4YhkL6pY5XXb0vOX87EVnaCjGPObFRXEqwFTpAcqiEVIHviufSjof
uQ+83qKmpyM6yJGdX9cXVh619OVZpx6HM+hgaHB9Gjb2RKGVfVaSTE5zrNFGnTI2wZt8mBYjUZ4K
ky0hp9xqYxtDoYx4gkeKsw8AUzheiQIT4l3zGknhkqJyVFAiM6XpnJfXMwhCIX8Qgh2pOic9CtBm
v5Xdqf2E0dWbv8rAqfmkx5Wdk63LSb8yQvN05i4bEeeoEqGfOBnzcTg8YO5csH92tDqcACliqgiU
v3Ft8e6dznCOQBQ694TCNGaauAY0DDvbl06fYPO6xUBFVj/TfH1n4CpgmV9Tg+2Cgk4oyzV/xUF9
RnmDHaJ9KhOVcYiIpnGTiO3JRrSZbWyyDiuplMcW32i35GDzM40EuRXARpjBJ2/+iPdkHvIFunoQ
sC/FW0N4Nn7yJ6+EZxis4+e2DOshHk7FM07xa3n56MpAO/NhHe9oE7RU+cmDVrWN/CBURQJeVTz7
APJtxDJdZYKpERZZcigAWAsqCluxL2GJu7OQ/5BO0FhKlcumPFQGEZH82lWpzGlT/Zb12Fiho+UO
t2OlTSl2IYI+rDNbjfANapHlO9IrD4A0XjRirYS4BSn8xTAI3AISgNlX3bbNL3EpN71chgtlQ0Et
l0kV5Dl6lM+WTSwKVpHvLFNvXeK0gNPU1lvPjWOJxH3szjzBHuYu0XwMk2EAqpvNZZbBpHWs5Pcp
9q+pC2eCNpSW0pWoZhpcclx0ZOUJZBXk9QgwMNUNg/ELx6+qfJKR/pow6c3cUfm6ilXbbiQIhu9N
VXm2IU6xEJJcd7EDi3nRdb3kPYlKrHFOxEdhizpS+FjRH1u6XgfuzKwVmoiBYxLL/QhFI78mVx5H
7qm0DccUWMp2XfTB+BJpMPiyYHJTwkgV/hSqnJ/OEl5jOvyRrehqsqLElluC8cDmFOwZw5xzlh1K
kmXJ8ltDklDQmYnu8OEkv5NYsjtNnebbvSf/JiUGFqeDAEcr9pC3oq8Aqa/o/i8GHE2aYHiiLk6m
nRopdbstYhR/Hx2bpKe59A4gCAY9RyBuq5heTkCUGbhDE0ugtd9m4gl/IpIVtP6MYum7YULyLQYM
ZXjr5VoAyzeqdiwFO4oLSF/wOuBQ78fPBT6uGUPw3weePyIPijBzxG40DeoVqjfc3//ilv94P4Wy
jfbbnlS+WTDM9yAksx1uda5ULYuXkcVyPH/6q0v4/eQLhjwArzyV3YVP0qg12mmqpYYAgjD1U63y
k7919btInx+hg7xbW6GqqCmML9qz7fC0pubtEOhTeJV7kRpvTV9vVZUs52lWH09qSW72lP5O0ga9
yPXfUpqewKCjC6wg0KhdJTd9E7vl61H3mq6dT8rMYQW8sBDl/JfNmqwqRRQN3IbNvlzDZ1xS2Bcp
LGfh0PzpgPTQRQy/XxBya++DnhuSpYD/nC/EJKN0xPoM5s0nt5ZUZWIuLVmeEQq7qW2ymyWYsDFG
1lJ+cZSFIIZtFjheM7yecRZ/J4kFISlWNBTr/V0PnWdM8FUSVMlm4G0UBudfniOhK4iTf0LYUfNC
0sOVzCulVaFfrB6Gj57SsjBOgH9L9l2uU9C8U1H4gk0csMGo0b7Ug7XRk/JANQ2ft0P4hLh+uD5u
O3JmG/nS01odWghhzJt9WcqWgEDuTYoGwzZ86BxhRBWP4M43x1YaYgJDyFVSbtwVLSiI31iOrDqq
Jll/pRNI/Jo6h9xaiY6iLlxXcsOH6EQX+E9RN0rzwXhF0iQb1Dxbnk1oLCy8kVt7kCYBsuuENWIL
4so0HUYMDwCQOZEmkoaHlOaI4ZiY9mRG3u2U1Ndwhak9QubkNnJs0SbHP5VYLmOEkia1fBAyd9C6
HPpe3DtmiM6whRNKqbyt7E1I5zb4W18mq/dmfpLSxf5toFB1vmnRd2Ua/lycrlrky9Oo18cfkLYK
lPeOIio3SEWhO7qRREHe2Me93wEzGxeenID3Q84fHU5ydV66UqNjCMJM22QDTKvdNJbJ1vE9HAPP
xHe9EymsoJhimDcA5oU3TyI+l6tnTjszen0VNqkpFvA/2lBfAlbSLkSeYxIVEALE2RcmOLcBOn6r
1XEV2LXIWLhRy4wo6lxD6F3CG0JxYCXdgGLnM1LWzCozo3VZ39K4HHsJQiBStDlWTh900OFURi4w
3Ry55p4/wmI2HraYEGSsNoxYms0N41+Vt+TByO5Ws3czsxZzO5bNmALqrhGSitZmM+5PHKKrSedC
6M/MsIRGaXneynTvvTIf7BMlEVAoTF3+wI4ncP8PDQyP2OX5Fe8bNAegt5vjRYk3xdQIELe7rT45
NH4N1cxvHPWErKJZ48NwUdd0dii6+OoJIYxDxSyXF8Zyj5/AuoKCnguwYF2h62SYE5slNGyAQDL7
exNRzaQPWUaAh0Ci1dYJLU4om22P2BMNrvmwMwVJK3nGQ5QiDiiz9EwttxUxq5bZUUIKowhTLFdi
c7qdlbw+zu/CH6PlyI/WKIICqWAMF813E5GL8yIp47a63akqMLx971XMrjHILeUE8AV13cVN9YzR
rGS8i9AovAYZ3R0MnAQx/RXdL5dR8v4piAzfSQFV+Ap8OZAvzvVvMIEysB+hWeoGZtwHBFhd77w1
crOvtJd7/O5s1uPT1WC7e9wOR0gEABqmd60BIEsrGGo6FW70S+nnndBIXAUHDJQt51L2ypt+UIZk
WFroaSsOHH9VPETAJM47SpHU0JOVU0oWmzAzrIu0+wAdLD9Yx4pPZii4O5AKdL3qQ3JMTkl0bqjg
D7vhDk6kpgsrxuruPfoeV0sDrYEauzlH0Vv1ybzVD+Uvi647THGaybNzRqWzdks9CFqBZYLgrrxR
vmFPEhQM1tLcntrL+s8NOE7kT7MrLKnDnvE+7Gv9cq6TRgs82kFnfzQP/UrGrM/Yyh0NhwknkR/B
9udYpymbcR41wUY1gnuLwPTup8zyfchfDs6oUHt8z7xqh058A/8i4+FeDW4jcQ3EEH3a7qeEUiIq
NnHXyo9657d6VV7rAKgWG68cbVVfmoPqNrJ9pObUaX38TYgxnCgw/rA4lraqeqqQ5ZchBmCJIDDh
aYGmGsve+JU6aL0ugbROlWPuLc+QZtYv3f9GHqPq3OuVqE/HcgsObfV/iSjiCouMkVfVp72p8o7g
4TDjVGpchiBzRusy6138ZwQVddaVDpMzWBuWzoy88h8biZtMpXoaaxvHrGnudbxCwbXQYpoalUDW
6qapDydou18tEa47CJJld1cR7EypuSZ89dq6vm9av1o+BIJEcwA643299h5GUKbce2bpN8itR9iY
9lJ9qi9lXV2QkWspZUyfZ2TQmyKSGs7iCfETVI96i83QuaRRao8m/QUEWU09ej6IkxNOT5DdWSxu
F/PzDa2KCx8PRl2xYrCvIRiJP1kOYnoRgUf6WlcCcxg54Gbx5A6Xm+LXiPepc4Y8Pe5uqgQDUp0o
av6aGpyrILgSBjmUxWbcp45nEXGKR8fpeU6IRnEDK8NanDov1d7DiAg7FB422JMHj/07ITpcsA6+
spTOq1biPEZbJsQeyvNJXQRFLG8ski48ct6iDemQ1TAnG2QYfth2k6nvqqJYBqZbeLIYYCLWELKy
W03C6nQ6wOoyC8XhTc4IIl+StoFz/iU8LAZ4+tUwcQICzLGCUkYDiLq+xJwMVzbOYThtc9qjCy41
esjDlh/3tJ591ELv9ncaevo+YCLTqIU3eNFWxJHcmOPxALAXxj7YFnki0LBLj75r3gxxwK+qh4Ja
lG0RAuYVyAqERBPWHQ44ssQNYIH3gRX9IItZ4xjRQ4f4Vu5OLw8Ysb4NxjrGMIAMFbdlWXESm4hC
LH5HvYswG3matC2TaCdMNVZ5R4aTX7v5x5WfPBIi3ug1/nbO3yt9qg+MdohR6Mwo+SiYxqQ6/Xwy
ayRLzmtJwun59ItaA2Hc9rnkk8BVVSKi9TFfoSwDVDj1V3OkN5RbZC32TfsdCC60BxS6UK3I3IAj
OHJLVCtFnaSorOuHhN+NsedQBugVELlJI0hwkhTKpqlvjoW1ukgK5URuimZUYS4GziswSgtzYvai
HqppcdDCotNumtxjPnYPzkmpLrpDLCEbBIhUgAKz/eJn0ZSClHFuUjAk+P2a/JnNCOskATFbq67d
/ocAzHJvmu03L9cFnS/9Rcio70WbtZ4L44Jv0VZnuRfvn9Au/47j3uR77EdW66ABW51igo0RtONR
lY5JuJk+6BXFCkjR8dss3KQVxCdyP01Z0WHKT8IVmbxsdOR58DM/hOnGUoPLBOSdOBfwsDA2bPFq
7AhZSZiUTgak4dm43jswjUqB9JVaulR4vz6zCMgahyfl3J74EMrkgIGyjbRbcMO339Qm3PqcCn87
V71uc7WLVFZi754XgMgKTXdVp7nReFT2K5bUxYUVDVUPX+o2Z+C7RgAvHYmfKZfLOkgs/9nVSCZ4
YozAvNR2YOTVPIQjiBI9cAGEqWNgQSXLgayT5LRrRbGuL8fz4ECHFlRReUaWCA5Fhr9L26+NWjtA
F+6iEc1/MFUg4tsFi9B8VdEeM6hBpmjchGFGYtxOlsCFQk/JQnitoHpF0ILINV8pzIqzp9g8h7ZO
CDAx/L2jpo7/cSTuHNmqj4jIvV8g5exWYyVTgwRrL81U0IjFFG3/q+ueKNZBWVRrnxXxFBLd9xaf
x6+Y4V5grHx3nkIRbO+F09bGJ8twH5VUv/Gr0W1WwUtinwgtGOEkJJQ94OYYrLItOKf48O9INKw4
INfPXFFgBTi1NfGTOHAZnKo2+LjkjPhWqoVyFibd2kIWQHJG/Y0vUxLW/oLUYbF14OjL0iwSP+jA
Nh+97okM0YvY2XrXN7ym6oFwlyIYNjdTrQc2HLGNvgrUqeo1fgOzYjwVQdyFNM9uozbv4iWv4P9V
C1JNw2skcTkcVWPlHCaSMY5bKtD3ECDOFKfV/DYlh3GiGs7mIoPeQvIq0ZFz1v8dlTYOtpYxemqh
lDgCjlH0aw2B5kOxGzBMXeOKNRZ1ciAmmd8QP3ozt0Z6/YIQtnH+yHGMTpyv71xO+fW6So9xLxO4
oPvYhnHNmKYLODlst26VpJkdyrtZTC+Nq3jaf/wD8Bt3vw2Sn3BiXWl20iDGx7pNfvO+Q+MUkpYZ
hxCcBvQtLHtgwG+JLc46cDFxci4YljqQqJBcaoAEwTzlFcUgbHbRiFF1bYYztAssaKpo7hpPqVMX
YI7hHpNnf7NmxIX5fSppnWi6lgrAF3EKzNLYxVYvxFOM5eZ2qzf1Xh9WJyEOjsrDJPgwhwQt0BAp
vVCNmWttZPCKhluzUZ6Ca8m/VtD/CZ6nhTz4ud+aiNqjpkgJ4FxkUJMM0LwV58krvXdkWUgZdaD8
tCmjjkGOS3k2s6+Jm5qkiaBX28mOOeAKjYaqIbbD+FUDEuLJCj9pHkGs1qLBtwLdsTS0GfVpORp+
LjXjViJrKQ186tCkLwB8++wHJkCqmu3gnBFi9a/hNj9xJk/oTHji7vbrC0ozxstE7iHN7bjJ++Mn
W6qX9VsFN7W/ufE0LBaCgVRLHk+UBgvV1E58f1whrqmzVJu7naWWwYWHqSgaRWUbvEWL570jlr5a
5LmKiFRcN9npbGb86cQMVlBlR5mKySifxdEoRaksvGDxO7UYxJBEJvKwZI7dAcV+0aNPCplHers+
CjM/CMqDwmHkh7ws2EfaOS0gwLKiRYOGE/Z2n945E+gkCOYvV2fo2sPQuKO7POWWvrd0zney48bq
eL9FzkQmHIz3oSSuAWxz4b55OUhbQmv+1h1kMkxJaOq6b+Gg/kHz0Mw3OK2O9JBkgMNWY/3ZIuTV
esCbaicX3ksDBi2MuhtERYXSdYbfhKIs3zZ9l7Ps7VMazAczSi7znQiBR5i/I8enkILVWKZC3wVr
CmwcJSEdC19+Knw4O05LimA+9VkGuQtpXC2Jj9IpF04Rz2cqt7LbTo25K8oHrc0mljr4l8ZL9lVW
1KWEY6g4AxYJvnbIERbYoRyXR6GlpPr9eK15gde7P7Dm8nrdqXQgv3Y7RAi4Kf0KircEqGsJeQxI
UHuluZWEeBtqFBbognghltCdAXemNs29kimwizs4YsRzRr0rzOgcVVu0BBQKVxnCta7GQhJqDED/
ZYQav9LVC08fw74U/tJxY/8qOcp4ujsYd6BJJSeQO2pyXeyxYPGA+Nz+0He9VWrgjnMeYxZYX3sg
CJkQv/oYCaK4QKtH5whEc2HV+0CBBgbT1fvJV57Q3AXN0IeAQnjFRP6X9qRfpO1kN6eY93H6LM7x
Aj+eBkYrSoOi3HLSic2K3B7jW3G3GNVXjWTdlqGA9udnSJMN8GDk3SQpGUrHZeoqqCuU/WAwWi6I
pWpyKJUOVjNOn8PtBciM6Wr06CnQ7W7ZYa8RduiraJPrCkDBnk1ksHK7iVwZolS3xY0OWh43Hkvi
brLQmUpKxmVyJ9P44YvJxPW65Vseb4rq2Myt0FdyqI+ZcqeyMdWC+WhacMuIVPwqUVAHyKKNrCb1
j5GgMn/fY+B+v6OmvLiGPb1VL17HFugxa1kmVZjpq1CQc6aHUZrkDfH7RUIaKiRlgzatevZ8ji2S
fAWIegUKMQMZkYUbcnO5Ur4CGVvMhJODVoug4vxomeosX/Vjhc+MB1mNP5Ka1kNe6itQXNH3e21u
fWui9y/DlaAcp350OB42GTsqq/aRQTUwxBJRCY1o7hkZwa728rHReqKA5VevjCti+Ju09AcLS3IL
9zGsYrqDHkYzZvFh8rff8Zuh40AflqqspAbvzwT/AxdFKYOu8I1jJiKSWZuQYN9ft8onSmMMgwFK
x1zREVaWZzP1JwPFwccLDhAlUfQVjD5crp7mPtySaANes1GaZFTM42R2TxjC8sadjxVvXkKw64yx
/oa/iddJPRWzTpfLKXUfM/kL2DAHxlcewRg7vHGSCqBW6ZSFxVqeolUU+Xmxfuv8NjvPeTQmoDs+
QQJ9k4l7oJ0Ef01HcNghD/pl4ztwOPIsQ6tIWUBpyI7CF7iWLgqXGsoPQ4A67zO2bEOaJN/yNPo9
nxleZIvq+aLoQUPfMnejd6M+/iDjhU7p772DwlW2qiUudwQ6B0tf7K/G5w1ypr1x/g3hY32F9tYO
ju1FDAeAIDT2l6U0cLRs5ZeWt4nrUty8bDlOrN7nTb7dpHlIgswJYruFmjsF6x2uJsWxw7TUSVOY
NbICeLiWfENVvyJgIyqhaHq8j/26BhbdDBF04NZ/6QbgYxJEHOdVAvEvPEm6bqiqMnZbGiKQE67D
6GjXG0661JKvYjwS/Q7EbXqbRJMuq6qvJ1i3aqV0B5TNYe8jPu2Jkwo9vCGOkc6y7+QnLCaCk5sh
5ZmNGFw10W7rDCkZeLU1M8Sxfqzoy4exxAoBVHBOLFhjPWqoh/Z8FxmkiLEAZ2y+8vN77Jev9R0U
j9rPonmQOLy5358YnDLzD/V7iwzDrp8T+ASavZpdx0pbkqfXis6F24P/lOZEMKmaXqKIgCsYHoet
G7/EHvm7M8r9KDI8OxXqATsMMT2S7oIR7CY1v5cLtxnvty6/2HpHLYEjfjFJ8StvOYMwyEJDsCdt
JmssaH+AM7Rwl7nJoOku5tydmTwHc3MzT8SNx+SWEhEIAIBNLXO/VIPY8ikCssqqSCEoo8RP696k
xgwsa6W+AbSQFfUbZ4e6/2zxoqGNkM5kswQa6Wt+O1PnmByWlFg9LPGazhzvx2pLfktl/ZQWAK8J
gDYTglrGsOTNOHw/JR+9Nh5EYZbSAfuVvINLbQ2VUxqKVON3Z0MLirVhprDvFcKP+SedRCutHN9l
kcDi/1Frro8PV41HZFWD+Aq9dXzJDxumEQ22m0lXPhi35Xg+8Kiyi217UlX+Z6vbixJIHirMPH1g
Wm8y0lylnyAlftoOP0poTfEPQ/CdR/oDS5NIjNo5FXBUSObsdfL2pfMLB3h6x7G4AIiAKee6ytJ0
MZhZ5lYc4F9uKQ6l6HY9Hsc6vdET4neP7hLyT5qZkOXqwPVtAoYOChuIC0bgHgUtxupi4pN5nvHP
pnSTqaNoze1aVUqWWuiZt8OGV3090UQrwCG5O2AoNRegS6o6wba+OrTbwoU2imotRp3Uq+3siycC
/DolP+7aINTU4Zclze+2NaNCg+0+XvNTAWivjhdkUcaQo4DE4/R5qVq5ks5Ripka+ylahHwO6uHn
ag5S6YpyNvYGMA4L3CBXLbHttaiFIpPI+Qgb3y2E6z/z6B355mBju9EEUrEWm8W2iJ4T6jFlaUTe
fSw4L257BAnesdDPBffPwbc/WZ4I7wg+p4ujU65//1Hs6AEcNeb+MFlGP6TFrEWckXSvlf5UHKvV
nzb+FgcNybFBYZPIDkDFVHk4Q/MsUIbJ9C12BV6+C18oKh8qq55MzHeuNsyP6w1jmyH54n/xIRaX
FoIVJGH0IYVgBqxWVOSg/fpf03sVES2CkkkK3wKsjouwv4H7zMeH810fv6PR76mv07BOAAEcVR4M
T5ClZffl/bN1/0XoFf6EacC0dD/iIsuq1lSwQ4adnIMI6o+Km2+GBDlTeIhe3gtA8BvdAj0h7Btp
+isx+qeY1Ox9h8C2fU/qvcMyQnDkK1pefuo2bfjBGEM7zuM8C3q96XfHkG5dCt31Fu0hc0Mho4S9
1jYIws2fNthGuU93Gy7rYqExzDTpfcW9lm6fJJ44PaEARkNxkLXxAprmfkSPB6afLXYZow5vOD+Z
7seXjTQ68meyhvxlUHaKpiCbtsOBaQBp9vOxlOTTNrGOpoQEbjdupf77ezD88tUYWviVdN8DbeIS
UQj6hO+vRv+SAFssBAvH+gaS4yKSYApM3FDP4OYabZFtncFAoz0I/akfo0LeM0QK44vf/VbO8Je2
frDH9mxFv/zUYAoB4qUo9aaCflhy4kQ0S0/TK8T6DhDAhG1CBJ3ugL9v2PIqc/AZgmrN4YKsYLaB
KaRqGmmACeuSG2aV3AVTgcQ4cPmbreqFwy8UDsMIJ5sb6PfuZArpaYMigObN5A/KIlBin3WWFmgl
NzuTxEYtj8Nnjzan+GgI+E+EGuI5d2/sgLryY/E2IThbFpYlUsrE1JwJQSvxjTmbjtaq66DX40y7
kzXe81OCCgsTsF+fTWwGN6v+I/fyDaU/1NdVYdCUswtFLAme/dCam+MOpeUt68feiRYXa55DbP0c
M3S+/ayYtsjGU0QqlsLdRqsgGwqOsuGUndDRMvmv6s88vMRZ+J+g5ZUt/+1Binn91JXfdY+he2al
vUnNVk+Pp6bueWQ+oUHC/ZC+HDnYm17IUlrOLZoGVrl301NPHxmJ3oqOrfCp5ibJP/7l5nBUQipb
7DlKd0eQySH+sFFhyOup1m+G1zUK5r+Cpv4C3m9L+sPV3apZmSTz/wupNRk0Kqz4aBXXKven/9ql
a4tClOAO19HRwPN8kloxQJIMMBY90BQFqVBRIKMOyNCUFIzIu/XTDNBMSKpBHsE5ydjoUFZVQxEr
QXAxw/yx5BgnRWU4WRzNWV3x/z1/fd8aeh9xKj7evSn6jEWGgx9BrLH5zQOfRePeUGXXQgTlzqBf
boGgSr5g1SByaGx1kRxApjPZgsZr6IWRw9gNJBrVUpsHupUB58Ctxozrv5P45BOkwC4GfvTOgGRh
s0RjV3YsRpB+Vi1Ax51gGJG99nIDlEHXb/UiIR43fO2/3v9TvdOLFC6JnDdzSL9Pe1kM6mCSeLf+
Ar/OrveV+kdEPYme/+OKAKr92BEr6Byx3pqjGHKONsAw2VNGA01v4DuyVSQDdXx0Gxn5GPcgSDwm
pBS5TrUv2llohgL4cED3AmB2cZJzyTheOL8O7CjXYZb8Pe+RkT1c+RFX27MoF9Y2rC0qcNjhrJ6c
jlrUg8LnJTORRjnWoBbR+J1sp8iQIBOLDqOs6HzAMD+SfqgDcXQg5bKVdvRLP0IOOsE74hkphz88
ZI/9uuJ7aj4xkvxsaT5ANaiAukJsOmXcc+YF0cBLZN8/IBvWlwHOnyPsE3k79HJYNE59lwCXmeJV
J/e0QDMV3P7YMxl2TiYFhdjQeOkPVGRePu4cV+bJK1x6H5dRmKvHZtKI5+9ocAlRz3sjlm/TDZ1B
S++Ip/lyEbv8jIWRzjiuShFxraUBwPBeIpN8o4cHW/eaTrED20I04WWBcTYJnyhnLlYjFd7ruhib
dK0XH/MqOHfmU3sE8yCjJSwomtMDWm4/VvRfvYEL8oyeWZIu7X3b/dvMo7d82Bsp3s1PdVkOLn5i
ntE7nigIXzQrZdFmU+XKiZsSBzdfPd/VXlvYd0WjkHH6nBABzHRNXRxyLOSx5tKN4SdIN6nHVwZK
kcTMeiGmBTYI9GkZZh9cLlHWiyc2DFZ2Jo3WlgaU6sLoRMYNJQ9fmZYcfWwR6aNctEpayiX47vYh
4ugnLHykDzBzkDUBya8HF4iYyTBUs7yT/pNSx6lXUkafDRXgJZzc9mLnumXD8/4oTGMpGduhiEg1
lpxTtCNi1KKZO8KjG0qwazS1EfQYZKUTIhoFUAb7z57zMU0n367G/wLvQn2HFjAkALZBcCEbKKKh
53wvpAK1iO/zj2ZMHC5Smo54a3gSyRWt6wr3abdETZmIvpqL75VkFtkgjSmAtlXTxzp3FahTaGDQ
tSMVZ8R0sUDbC2j9CbNpI7ShqQPJUx8Gz/bW0A/QgbvmppbbYoyvKJDPgH+alKtubS5MVNLEYt46
LHhxNIg21ICd3iyWeMJ8sh3fjdydpeiI4dA+QZ70ksNUGSnnM1hXQ/BqDuEKNQ1xXGCr+z6Qcgi/
jy9RIkAeggSR6ZnWEaFSCoOX21dmosofD80TjNf5SDDF6eSe3+7P2eC0150Km2GFCExynXeex4wb
lyVrcsOVTaTtjUwhX3EpIxA9q01x15xSeIgfyuB3THtxCgmekCzXV/BkoOH9vvP9Cd8HZvJ2UK/V
Rqfkwg+lwq4lckosBePbRskptH5THGV/EYXubPNpNwOxmn4qAd3fRiNSg+uh6ndVjzBZ8TPqZCCS
308+ML123z2QJPm//I0HVAvfF5l1/93jFzl3xkUQW1tNw8zhDfah7zrXQDklfIbvhQuM3Sm5HVss
FPNwlHqFvotpsilklWvpJopvd76fCpSrxDUGUoeY74xAAGMZzFQ/kUXesPIh+B5S4rF0aegIOba2
HIIfLjTe617LeRWQ0+fuTekgm6T6+GGmBxoOGn9fWJcqs62T88Nfw+kWzgP/hdYKkx3ogxBgmC+2
/OaKbc3ShEMwM07qiGEmvTVRJ8FZYQCfNTJhRXu7/ZKZWrnb4+BvZQENZT1qey0UCPy1TDapvDoe
DvuzSAzTcd7MuCQE+56GaSgPLOE26XZ1UNjHp304MOwX6aF/AaKdhG6urcj4Rvn7Mb8i9XZ3aC49
+lynsgHgJkfE0Bgu3eKJH7MBBDA4l6U0AntEIToQOmTv5vcGvP5TksbwUgZtAo1fCjvWIQrmsz9M
YSeoupBK0xNxsxJmOdjEUfzngk7hZ6LQnTF35y2DrsKkUNCBixsso27zhRURT03laVX2eb37BziE
SrPJiGY0qVF5NNrW/5WhejA8ZXAgDz57BhItgsntLZsdMrTkidXgx+nBGamAZEWS3bKeT0c2sHpj
aMD+RjVrtHeskn7MqixkkAe75R+d7oa2laAhpFq7/9x1Z6cEXoV7PxhxnfsqX4JzxgKDdMEE/yvA
eQ8qshZJ95KZ5lylWeJM+TLgspLrm7KeqrnrCgY/9j9GQlwQdUW5pfhKBweZ8388B1SdMtFFHbJe
O+7blbiODOp6GUwnx1hh6XCrbFZxwmWWtcyot3g0o6thOjXst8+aM4gm7u/I5qyQbKzu6lYoE+Tz
JjalOLhGf/SLYkhdre4WB/Qp1/OJI3C2muDXBkRNeb2/nK3dBFO2SCKRa15vK9/PfCWZR/g9z2i0
KQHwS0K67i2a43coasa985HgWp7mOh4rL0F8XTYm1ICLgc+1kUr8dhkomz4j4YHzN3lTpqTzLtIw
VTCNu0VbqhfRNarLZzgbVaOAHPLqXz3z+lF4UMe8fcRB6WGlGtUJcOqwOEemA/PCBKm3LTNwDmzz
jW9MncTQ9XBTOUiyAK7hp3EZJGouCgUudsWuEuJsOzTLEBa3FjQf4u2ohN/DSLjElX1KGeowQXuJ
ebSJ87rTgwMuIP/cmsovKV8WfUHDNmTdNKRVN5VzzWbN6c7Knw93AC84d4eCUJvhDtjpYkOcXlRf
m3vXjMsRKZtiyh/RWicCS7Bz+sehI7ZiybX2Qm+6sZeDyszNNcvHbKNljR4USqS4DRkPKQeOOHlt
70r1pkBbw0+pp8dgb9QOFJHVadNT2sVO+UE2R9lqBJqWecOBzKCHZ5Wb6F1W9b69H+B45jEXf5Kd
HiFm0z1L0BhicHkRnPcB7/fPD4UxuCRSnDoB3OgPu49kr4UU0Vt9uUtZUVAWyAlGa8SRRAzscRpZ
GNEOW4dH/yXFFkoqPtoWOaxI3Kxc5EA+JekQifArKx+fw+IjEYMyvRw+B1LOC6hP3nXKwL9BD1Qe
W4lmmKs6zBNrEsxtBo/gGczNh80yUbsvTXi5+cAPJ6xwXt1UxcjWeL9Q8Ve0sRLKMRHuLE6v1jxX
o0B46GGA7j16XYUKHyxs97OOC2ojsimSgyvBI8BV3O18Sun6myFly8/4iuLsKkXHkw5zoC9ANQ71
IVQR9EdjyA3SdEzjT8Y6oCxVG29B6/emw6TOmwe+sN5gnRQJSIqYxEqR8FyWNnEDGoBoaljchSqa
VanbtsTll+LFVcCtbHi/DVvHHFFQX2vkoxSUk1iR1pwyMvGZZLcI/aQ60BaqQSslLoFdWJaWh2RS
UlgRSSfgIxCMc7Z/33MFxoDtmw4NcDPSEeZJ2hpjEK+6Rytl9INiF/P9Js9Jpmx6zVDZWmrNZ5CB
0VSANv9DenLlQQJ+Cbr9YLUDRtL/L7LIFVO4RkohvaXS1IaC0p6tdMrVbIN4wjkiFSZGJafGpf3i
DdKtJ/aUwz4nsu+EV3cD3ALimhvj8qUA6EvhbzGBIytK8orJku/ku1pT7pEfn3wtB8R7hpy0pw2m
hRdDr2GZZ0DNDlcIv+6dyghI2TZbZPXPjaJaCI/LfnWlus6CtmJgc/uEAXuDQHDc2SmZi2Yhk/y7
2ca2fsbmbe6a857ZqyeVTVokH01aY+sITLAyLfdVwH+jXqb8vcIXk+ujHybT0kzTKNut4l1GYYF5
2Y4UFxHRggySuEHnAmLqkpINNRC6HgpICs3S7RBcd0BgUpaQvzwTHDATcBcAmE49gj/mta+lG9pX
kHGEHOreScEKQgD6ELiV7HBmLQe2LAjJtDEx45FFaUyWSTPR/jzYw8mUeXI/Ps4ycmyrQ04e2aNn
cQGX9l/1r+L4PRalfn9i/QP0aqQecPr2xXz7Eg+1rTtLFgRT1JaVclGvDsgMMZFN3nBQ+qe2U5Bs
vFrZYKHnKxqNsxUY3n7EvSHrKxy9R4/uuppA4qJaJZxMIJVG0MlkjSvf5DIJY4HlY7uQ0aQwG+vb
1bYHk1EkaiKWkEFGz4il928hQQFbDq6r2S6Srthl8fk0N4YS2nsKsLopgGvRDQuxCEG329cgsJzL
8KbEmj0eRHGAXZfhFYBC2kDH2V3u6OvHDfk830wor6lY/OWKHhuqJqmLfvaW+Ki9KJu/e9zpQqmA
UGOPwNC3rgJHPIXAJjgZzTQiPC17eA48d1E9yma4LFg5KCbF3gNRH1kSEdL+rrk5a6XLeD8gk+hQ
p+eZR5AqTa+vroZ66tiqvGkeQMKIoK7M2FJbFDfAXmJYETV63x+T9O6mlfM8ePEb0/70Pqz97f+v
eS67vXfgoIT7NrsUH8lzeX03eaaNJm1IWA4BK4QoAq+9xmlLn2syGkh5T+vMcSQ/stnbF+Yglkzs
lU7x7XzU/3r0HOufSMjml2/WTEE7kdo6BOGi+Kw4kq31vM9s7EHKeNeXBf3f6lNKSz/e/yhkqXJt
bDXoPOQQM1wg5Sq9YlyjGLPZT2x2uVnSHCTLcV20+VneLH28kBaoF/Aop6if8yQWUQKTVYcEEHxT
I8asHyOkCinXBkAa1ctjYZA6UaIR18v7Rt/F9mrxmDKIQ2SPQbQAKyyC3vG/Rg3HeUKv/iQg/K05
JX0i4T1TohQs6qGv/ZNYI9sj1T0hFi1BgDrQQA6rJ7JIJTg8bsRdnhS6xTsuEukxZTibJ1sPDl3M
FZNxGeJ5gFNROWVCMsO8tPHsPDXHxOPJ3/6YV1KMq9pmRFGe7RH4yo2Tl2vcScbEtq5i6ZGtXPyT
MTO0O/JmL/XR1dgnKYd+4ZNvqPUb0t8J/ReyNUDl01Z0BxKBCgSiM/rOS4FIwDBcLQf0PIHmSzC1
H7wVew3ChHUb73Txs/n0lD6yhZmEAssqeChtGedh05Y7QpACQV1r17Y5h17dY6oQFXfpu3XmYIfv
wHFvdrR6GQDzMkY3xup62Asyu0pJUNDhRBsnoUxfJ/HM8qxkS1832C1qDcN5nDcH3X+bexEf/iAr
qyrQMWarZx6HGbbK9DiawavX1KLKeEeXJc0hvaHUf2wDPCUaWStaUREfCNUdI6Cr5FUgK/m+5jaR
eQs2GvQUoal+/vpVaEl4tUNdFP22eYp3JtdUsp/h3ocYlhDzE27KibXE8H3Y8wpfTbccM7bW74Ve
Ugq0WbpLMa2ZgvEcybMX24bV/nqz7e25eCfSnbrc52cdZX1EYGRK61C1UF5xN6GvsK4ShRE1kOf1
KbUOtty4XYt2jDEsy+KkNoxRiyxC7iU+m0gn7fRwgtihSFRtOMkRJzDb6I/i7hzdBKPxjEnmVSFn
+klyIt2nGMDW5cT7yT5jPY8otDCb1W+8x5n5hcJkrUzNR4zHBHiFoLu6ZGuyCXAfAoYzWrAYjFDG
i/YKQ7z3g1LybT5w7yNZQhFi/OCxgZVRRoLYaX8vJgxhQHi5X5835MZl/H1hgndRx8b07irwr9DA
15XD6hSfLiAabxCgFBUGFgrGkq+vzgcz0pz6xaxCbddwiNopgQ74Hhg8Ha9YuZcXWivauQ0WJXmK
uXFqch5jzzgLzwWcXhTC1G79R4PVsRwQhD3ND+A26GvSOfTNUs17wKuqjyRg3w/3XhNwGslI9UHd
0L8aL64D0nEDGaDv9yAt2nsA2lF/ylIixKCXffr9nVXXi9ozweWrnpM2cnV3tu3aGAn7GBDe/uYt
oPgu7uIdQmJ1waDjn1yrPRpaERxie9ipBKPn52s0YvaVfwTehapeqi33XaVMXZ+3kql3zy2XZVyC
rGNDVN2YWjqhlpiSMhvzO4KWnjUscQ+jFtk7BCITSAkj+VXIdYwFF2PnupKgOm95TQkXy7cEdTfX
fwTIYMngT/02cqB7qm17VK8ZFteqqesQJiE6ZJzc1mMUdsqOetpftzka2DLp5baGxATU9tQmT4ez
H6ZXYtjX0zIpcuOvsSUqExGU/kk4nU5Q5NSxT8VAzIcJIajZYxUJMNNfEu9Nva16HNcNW78moQt2
UpzGZhwRoDIT0QFL3c6bMPRuWa17fyagb9v0f68SsY5WCxIqFbdWZvsyQjabm4vgJ2PbebG2DbMz
e86eO6A8tx3LJuERs0dDYmJ6ilOOjqYZeqne3BPxshbyDQWhHhAKFW9SUDl9FpAlWK3PP6B3BOpZ
SoYsCLhBdWrm8zkNk0wDYBK68O8G2jRKv4ygUD0/71Pk9Cbjmr2OxWzuD/ReXabfJNCB2ODR6Ngg
hIkzZ9mYAcFZ/Jjics2bEizVQvCLJPtMwD8MRTnXdgNZHdeDbMdkPy8QEwtUgCssHML8Pnf6uS0w
Rz3nHv6mznzC0oWC2Fq0sWJzSAzWovW9qVH7UDOzsIJAuOF1XarOKW88Xa9/cgT3TAiVw/lI2a1q
PmgrW853OvfYhcZBtwlkQ+NJOtZkWDeM2ToJubpb/BmZfE9cAxxgd91NiVaXuNOnz6ohkgkY+mWS
pGGpT2KXrLjiQw5yf3kf9xz7bCIuo6R5PDCodhBMVQxeLlCaXzzpLvzqPVGNMFrhWjT8rEhMS7N4
Hnxjdxzo7Hs3IrjD1tPmZcK42xw022JB8F+pqeHzKERG9YUx8R5sqXanO83KlrBzOqnEA74ymFC0
ICKYcAE+lqQla7AFbwT/k6fS2HKZWh3ieG8yEnp+KOhNx0ml2mv+KIjmS+Y6kUxSCLWNmJpZyZMm
Wt9O5vYuumywsGBl6VLegBDkrXDvg69WmR4QaaObr1DHup9eoMY2UlNuFujcJSyxo3Xa8MHcC060
WH/UD0hLucbJ9jl7F9MnFEgugjCV3nGNZpX+xkYUwaMo6iSEzAzVzbNnFIho/9ExmgZBTq9GZ/yF
uy/FpwnrCwftGJ/zCNiAq0QR1aHVZ0dGit9IiV/qc+m6rm9em6NyX6L9c5HJ7mYaiXeMS40tWWcy
twQR7lrlUYWXGFmxGhZlbHVqIRen90oaY+Q13Gky7/+RzioBwleH26nHLrRyeS1YLetbL1uKW+fy
leeqntEB4qxfbhFIiJXyleGTQQ4VNL2uG7Jmy6iZHabw0cqZmztrYVXyYSLCrkMti/Iz9pAqOX3m
kg6nZtIIzzonl7TM0Mv7XaUqkdXdgHh8PBqIIE90Xlt8TS8BupUTVL5whTShmWI5bWQkwzvZpzHD
b60ikUE1i+0Zota/XUi33lPmY0IVerE7DkkOe2TjVM6IiwBzzPVB2Wm9gk94g9LNf0zkjMVSGamr
RhmYfN45Ec1cxZ2tTVelQ622nf5ESPoty/60NsZoMOhrm0kXCL9EMxUdNfa7ma5g1qffUTz74vAx
h3A8JdVJwcioBkBVoIhwc8op5iZcweqvUlzEwwffCpF+4CEYq3ia2DQEw93xnWqYxCy7MlfLwuZP
y/sV+T4lvcMOknoG1RQvSs3ygjmo3k1V/2Ei6TUpkdVqZ0cC3KlQ1xDmBBOTmIBXl2068AbW5QK8
wabs+kVS7240zvo967WqXmPB8SwZdTzf5ddvyAUrl4savTBgFrWmwp1X/nzsQfOdR/bUf7UtLrfT
RXq2Kx/ZxCdm4K2/yKhlRs1ZvYzIy9MnmCDqDw4LOOfNTOjST7u+X7Xu9VegW41A7WyAZn5LApOp
fXdnAC4PdoaYK+MAq0a8nhwQnICeVMdAwO0FEbrn8P+EpAjmh2Im8pdyEQvZ4h5ZEzXX4qm3d9Lq
B8u6XqmB3hCY8yYMTDbSDNv2YF6ApOzEEzBxpIpWeIXLzsfgULHC3yfA7Qgfzpfo8gb3MgTzIbx3
K1W1DrhUP2L5g1jMcUfZE2T9kOkaDcH0bI4XdkirUEVzk07Hqt2OYWC3FwLLe2AHvawy7hUXR5Hv
vO4LI796GKl3T9mxK6TNNFuXVs98fgZX/lnfvzl04+DADmSwP9DSJnD+jpK3DHYfAe7V160F9qyn
uqtTI/e3J7Sd0TPx6WW4xIrJr8ruELpKtiqZSj088lbOojdN4i+B5OCblXk0jb8LSZhTeNZdFXNU
iliKqwjuLEN5RUbyHQwPImHhEtHwkpv06xR/aRkxJoteqXy/VOsZrEQVVWYb6ztyZbbk4NzTPnqS
2O+BxIj8a45hlqyr5/47gNh/92ZMEoZmiXU7tUxf2ZeAnCZ56ZOpwnvARJ1pOJBRQ3Rru4Ysrzpu
AcovL3qTtRhP95D98doU17ptvKX8ZgCMFUqXNjfWgvZhbLZqg3T8uHZ8I2JrlcdKntuolTr8KmVJ
dia4bLHIs1PcwbDkFwkduEx0pbMwE7dbGYgUZQ7ki3VAxwzywXb3PFn6TADvpWUwmfrJ0i1xMFAm
/IHroh2yamg5kM0hCrO6oEiQX3W6Aumf44wF3qsaTidklLN6rSOV6Wp8A3uJdFWInbCweTwnK4cI
ol9M4SZHt1Bep6J27D6QtEagPKz83Kjz4gpFc86SQ7gcY41IAL0nwNbDYhim10m003d7CA12PWM5
iXNFxvYN5b/vEfg71YK0h/2ev7VfFqpiTveY6lLNh0FuF5Ua3Q43A8CfuIbZb8fH90J064EoGyLz
Ys7ROdlgPOrR6maSp/LlNufEpwr1AvU6SrjUFCUgmr4PIaLTaDzcTbgQZykZAXQdOVQVjYkvghSz
Lptar2TZpDlqO2twDX/1WaB67bVri//jHijgvrqpy5foZWSnPcytf3JiPuZkbWNmV9tjQraWZQZc
dJVdnVDYKnzjCRWdQrVAaVA06KjUEbsGFPWjMX68LfLNQGqFVDI4PJz8Jd6pCn/JFCW+qstzOeFX
janmSqSlvq6u9T3roBBvvDPw8bbCoxG5AoWdpeQr5aXh21QmfsiUslwGVU+6DS0eqj2ZECYEiz5u
Us1RUFsauqeEIOls9NeN3QTHkFD/GDkjMGUWBQnNERbyhTXB6s76yjcyjhZLcVJvAs5vkEXXK1OF
AU8kHQ5fDB8xLd296RdqHOc5eTQ6a3O7n0JzhDZtz55/nMsRELLPa4dF7NUCDFPwsYhNk1/I6SYl
5JHkbvRBAzfM2B5RY3Gcz8pfLOLMzWovKteF9B7C382dpFX/glx/qNITV6/9v2pXvsVZxUAEZSkM
dpsHPKU7QSc80vBq8jBxMPP+251eW80/kz3JAd94uilMQjcUVHruMCDHu5IbuWfNDv1N4g5ATE7v
XlQlVzz8F2t0VPuG8NlXQcCKCd8+k53mBjjFDvcBTA1r/FouYGGKSfaKjm9pY+wKMl6cT/wjE6sJ
cpigmlk6B7giyNCXEs7NHPD+zv/O6dqkXmmpi2zBtFWiHoWVpqeY74pEVteKa10TOypp4XnZFBf+
rbhccEmIafeIViNiSn2tQKOHQ2F+K01mHa1/4LFD7AZ9GqcsrO1CP8+fzFQxUCAepkUZpbJkv/PN
9lnAP+k0Hdx6pBes9KesFAzJ7ux2dAA0ZKMXVayBfnbaLcoQOEn8jDEkHZZTU16IPF2HvptOij8E
CH8UIp38dSEoFkDEjZdrV+yEH6uqY8V+olI+3yoHuR5f4VZ+cDdhSU2SvV899cPgJAjJx6nOeOjJ
DDQQpLm4soiIlUzzq6N+SBheWjVFpJmniwptoth6to2+W9IqGTtkf38Go6jgUdRX5TsAdm8KZRsX
p1bLDJiChQzk4RfKFsQM8COUZ0+TyjlGXt/qJ90LBPS9uDWNeQAw/YuUm0R85i0cdjb49g61Y10L
9sZg0ey6KJ8aukon9SJ+KRkxzYQkW5UMQgO4KIKgqWzY/eU/Prqy5fEc70nSC1JoCo6KgyvizsTE
Xyj9c0KOq2i349uCHOnK/dR3z6nOTA44D73rNoyDYywjjt8tnHXmM/NyjiTjN6c2BLJ5X7hwo9nU
nF+iZaubvykHorW7bQfpsWHFDNeUxOR8si9ohVlHOBmOaQNd2NHgZHhBmE2PF0leMa6uIbA7u11v
Ee5NUACGqMilkILpF/e+LCyA5xUf8OqoT1P6+0s9bg9cxnWel05rir5xBssA+ENjD38HCyc7fkXv
XQiPolWi6WxMSKhpo8xeK5U4I3Pb/VVZXwUXX5FM/fet05moHGAQzcru5g5/ghMs8t7IOW6HfW+R
VQ8DcMGzQtLWRRF3kpPxM+916dhsLa0Ef3LtLENMh2iI1Q5yAqyVYtyODso98UFIljFNWkjmvu+D
GzNZb6nflSQAF68uuakRCUHboSKVDYuc7LXvtuH+j0xql4qfHCeP9D7EetT1XY+txtio16lBZKI1
qVLenUk565oJ6C/TOt4nJofh9io7JuRFACdSXWusb6EqG8HJaa9cOwtiewe3wzAhcTN3uFhDKZzi
4cmaPKN+fYM7B2zhq3piTIZim4TeCZ25HLMT7zRqGPdWKcOM5nNAxakF+G3RsmAGl5AiDtsrY5VZ
z9LtyaFUG3MZYQ+iBAA0jTS4ejswugYjDXz8PT3B7NqTbXcxFKVFhRew5T5wYO98PaXYZS0oTU7H
q9pjaA/qyxORaMG31jQju7i3f3287H2PnxOpj6RYyVkHkCO5pV7a8wfL8Y/yNabiDqRbl5a+9Xgd
9BRpP7YoQzOs3v7z9sx73vP8InHbNo6ANBJ0//iYsQtbqAr4GKkgYhGk/Nr2b0wLhuXyUWqyZkBs
xAYhaQ9n7hV6UNhx3K8wSzYtVa5iqYB6rEb8vxauAS1XlXDJAE2Tiam3uoVDzUd772dH1ax3HlnB
nHd4QnDzaGmpVYskYAwimxElXN7z/bj1o7rXLCfrzdPWCVVJO1sBkKgaZTHcUm9JcioySB+O1Uj2
2PS8mv4A2skPrQs1Mk/Hpnp33qOoMHaE9nxBKRL3ZG3Jdcu/iKcdek/BeX6AanrLisRaImsJlBXL
Bj2OZtQdvxUN1ceESpMcDTCNgUq9lvFvLOLagm+SEHW7FinyqM0p6XI5WckbBtUuz1TpSa/FbjoH
n3sulQMOTVAWpPjSI0SGpqGpWFojfsSrhegVU/S5lufC6vrL+7rP/UFM8dbdtrTWmnRaymop/DuO
7iHexy0uKFycmWGbH04cmSkeRwyyaXFGgxu4J0R82A3qvQVi9mubie4zxALCAZQNLGRPTd0WMu0Q
53Rq/JEKTaH+6rACQPM+jQXmynXXw8RvEOR4OWNrrK+0wAzSR8x8JU762oGu3NGcAGDNSeCBUdB9
m79KuG1dXmbOGDLDTxLOwyLZSOkc1qKa8cq2Qw7rLvZtXiBKvpBVpyEORXM/OYUx2IS+NDlvIs8I
SGdhlkW4Rs+sK+KS/4VFP7Zsvf5LxUFmUAJdeH9skGhSisdAjDAaW91HFPOq931KBAcid/XDi3ZP
s5JL0q3fKUfZdfcwYmwObXyaH82s1Gf2BBmVzGtR5HpP+XA0BtREsHMOrrqU+iGU2mppXS6cR8Se
LuQvKOz8fm5ogL4Bbf30UU3b9K4xHqwbzW+YtInrbnLJ2vJtdDGr/cYeeL6fLvXVBokehBhqXmUP
Sf77AymD9aqKBBeCqLZ2vk4aVmz6hgcLQgIF97MbW09k0Oa8y2XoIH/ax2T8KGvPro/P3Jm9n7o4
XAgVs/2JmrdJl2jjSm0HReRip1AOewmFGRb1b+4bM2plZruEKWHfw926oTE8so6p5AwpjpvmWX0W
yZBRJ/5fzdN+drLgT2OaVZrHq/AdeknyspwqMRvhTyZtxpW1rQkSlC+Lh7bl+GYHuemDqZmkf4h3
osLObTQxBXkC6dK0fq7ZQHcDPhONFY2YWqh6jxkLdHI6RfSFVkslMWEkl4R7vkPxG2UWsp5+ayiR
3P6leKrp20YrZYHdoSVpVTTZlnPwXq8wWPop86qoI7E/Zg/smYDdJeSrhpsYP648KnFWToyi3PcX
TTDjgBXqlN1+q+9bAfxJyakDGPqPROp/F3DsK+UUtgeNnJgRqgSR4RuKbMsRAyTbe7WZxNsrsen2
aP6maaY8pdgkLrtoTSbcVjF9XxUyD6y3bEv6kf9nVeraCUgUJhXYBCkcmmWZlRSDWqTDcXH6d4u1
2gHjgv+3t0mWnwh2fO3Wlr9+TH3O2IQHuZev9QzjmM68UejliQ/j0FQRNlKRmt28Q2r/N2vpzpVv
wqZ7ReluxhnPORizYeKwfi+nRb8w02Vsbx0bzSApQoRRkgVAoSVspQNFNF+BPWT00jixjF2BPGz0
NRbIbA7YSZ8QKlVjwunDDzmkk82FQLTkSAickw6gAolZwMT5ZR8OW4fmdf+ql6EUbhsHlKsvi7XJ
EbOLHnj2AIt+IjIfm4oxGrPdcLAAw5JsfTjCEKGqeuD4TqsrtYFxbV2FMSki7+ZJdYWJNYIpPtfr
kyrAmfpBDLR8sHK2WLfyL1bpDoNr/FPPq1By2nIgmZAyowASV739FONPRN85mWYFXMhZDEfdd2oX
kVWQMy21awDkfT2uTTG9F+P7VyIEyWhsDNvuJpVVIUTe8VYC//Bjvxr9ajNYgdElFgLjpyFjIOt4
YR0JTBbezy1FP4x05KZpeT7lTIMRnEdlddZM1x1loSP0tNL5NsuxTCOlOLEZvMfd2MmBB/gbjbvK
UOaMzy7cX9D/ZKBLHSrkMYkm8C1E7JbrLuydi4iZ6CQF7MIbYunPk1cWP/hd+9UZNJjsDyWAN9J5
chAS39S1JS/KlDUSZ1b5nTjN3ar146Em0Qxb1POymwg7m7Q0f135MTv9/N3ZTQkMdFZ8MU3RlQ6m
Ku90qkWXVbqHnBnn3IHoPG1dTD9MqjzzGc2xuNQGc5t7FVAX7NlL7ylW/SSHfEGsI6bwT+2SktaM
MemTjMmjqDhoJ9VgbOSqIvCs3urb+93w2sMc3vGySebRG9nZwZ6MR0nwAXrFhfFXY5ZhoUjL6rxn
mmy8MoPDuEHGVsAWVek8cBFOWssHT8OjSfxwqHnB9reDWh/RV6qWpq0CarIOPS93gKI21wAtdt5Q
drmcs3qQ8K0Kno67RZ6AMJ49xgvPZv1H+SjUiKB8awyEPv65zI1rOL2o500QsRp0WyYsmUaK7++9
zlvlq8o5XS5N5Vbk58Q2cr5XQEx6Ha2n5VQqsmStt6gD0RMTFixL61wZeBwBwmArCGeOX5a/6wRM
Us8m5RuHYXXG5vc7Bhef6f1h04UPJ30keF6FoF5s8q6xYaTXUmNZDlNCgDn6w0UupHovBElil/lV
gJjLT2clFP3DGx1CBQDiug12pESn50ROHh4b42T8AFqX9OiBwr1XNlBvRnnX2eZT3SsYyU5evdiA
FrYTOIHLXC1Z5RFZ4kY1zwDJ2s+nB9a2g70Pq1pS1PmZo7IQfGLwUJJ4EMvz7qRaj3sPmPIUf/XD
lyeI8QxZnbPtOoJAa7ekbH1TKZG3vAqKUWFDwfOZ3mR1Hcb+AyhwgXtgBRPRTRhX5fB/OoBMXB3y
ngV3mv20cjyt1TQPaVEWugKDizI6dln8Wv6/JlgCFy/8dUP1VYix+NGk2irNIZ8RxRanUIoyPP9y
HTQZOIpqF4D80S7CFaTUPKD7GjlxYxIVLe1G9UGUdvJ4+zoWij0RcH0W/KfpirB3kbvbLAY0seVl
TaGvE6dzbTNSJmVEO2QcxZ+k2C6DPMSzZO3lPm16JedS48ZliNktsU3eOfCLgww7pXVdGg1naDY5
Z2CZmAZR5dBaAgdxoJmPLIe9msQHPglOkrgtsPxiHWIKIBPW4Z/om0+D7scJI96t6qad7KbdsF+6
munemBj5/y9me+IASBX8j8PnEol7Qe43/HN65bgFbZj5fTUs2lCeIYmD6O7BYjspe/QIEhZ0IYwB
jfZ6vSsKh5mM14tiNe3EmxEAk1RER5kAZMntwQ3czJZncw+b1KOeEo78G+j8OXn0Iv3ohKDQm5FK
y78Ey4w5v0nOUy+yIGWWwmJ2i0Tbj1ZG6kn+FYyYgoRqit3J1ja/GVRDHmc7+Z8wqiGbH84tDs8N
jPlXg7KlhagDH7szfC1RmTGqj4dDnSUKMRRv8/7vkYyz3lsb4DyCi4MgXi+YULZP7gVIPGli98Fw
8H+qaoyOdv+Qp9WtQBY///vp+X9zcq3RjpONZwa1OX47d/GLhPdA8coug5WriKom5eOl87wbcWRq
WFFuno6MudmY9lzHkoEiarQwMgYlWDtq/yawGCpr8syWxrexr2aTwVoGJ3IJaSbsF+CKgkHmIFpD
EkgGYEPxA28R9mSLdL4NaFtEnV5aLreCvaEMapo+G8HTzR1jOED+J6RMdzODclz+kRtVhMCzCIMd
f53rdKdG4YbW7BWLPUtkZAQ0RpGFTOamMIn84vgAhYZCu+vHXarcIYYO8itub2vbFiEWQ814x9Ft
ubrIHK04oTdC1RhYM1p+cpPPcngEL5wnpQl1xVpNTPipI/FZX4JkY3+LFY9xJ0WSz8+QKAsAy/tr
QX17yXVbomv8Hq1RGxEH2NwEpP3kLxXtOFVbaYKc872Me5QnUj1eC6oZZPGPM/oilw5NHfi1l/t1
IGUKfE2/eEbmmAk0ZITp3k0lX+BosNnGqtuxxiiLiJwGdFmhyyX7sMFd3W2t9ITF/1ZepIXp/qqu
CePnkbGYZKGZU1/cstInAQ4jjjPF9GjWeRJQ4lPvt+disR10GlvIRYp5r7F4hO9NcFzlWfTqsN+x
2HAhkiONjr6EdjpScm9QySLS6g9eq7uTzpFyWViKf3LM0w3MIpuez0zDsbgrYmZqnypQp3uPBUK4
NcDW2ORBVf2BT8VU4vBKeAGg2vbgVNPV3YQ5oUf6ukiq+p3KfVMhEltsJOlx6EnKET+wucBOHzIF
51nc7RCNBzQjkg1A2ImaEpT9mS/2XYr7Tzv9AkAQsLcKSykW3x2Nkck0cHKUpdu085L3Yu1AWomN
6xz1hYPrYLQb6o3IrKImBt9FGc5yrg3BZw9My2MjWAwxAHjz90OLg5BTMageEYiSTDJ9Hpbi/sh9
QQtjmyPHxc5JJF6MIr4bq/BzpaUP5CLEystDHtVv68+zUoSBO81Q71peHhVRR/TaW/BXyxnerP2b
mM5DOjurXnbUF7dpcxtZR27ijxyhsSWYg8AxkdlnCvJeOwYS6sGlrnEkNF4q59v9f1eFBmE0Vl2v
WnXIYP8EeRWyeSE9bHFDxomz5TH4p7PEqCTAmIEaehGitfoUDoJBFMHX20llhD7daO2q0jjc9Tlf
l3y/RNdMiOwUrDLpRkKsNSwZMkGOpRY897HiMLmFdOynekkvVi8Qas9FJinmx24IfKvJKisV7Zjk
9IqakpW6UaxMJMFUMjH5TYB/W0F+UvOD4tZ4hXb0yitPV8lRqH+npFnS/Dsi//xTfqRyH8/rcRDo
fzSt/V5LVg4i7xdgNdrF8Mj1VgWDbHveXN97aIwEzehVc3SoshE9P6ABEsfrnXoqqsfIuoH1pVug
KyschrbCuBnxg368K5KvPchRu3t0/+Bgvfbyr83OK9+culIjVdeomizikrTXVoSARIgi3XngqZpX
sWtuHyBVI4HS+EFB4Pf0d+9vTPNmoD4yW7S/jEotJlKsUNn9bAuAG82z3LTKKQ4VsI+jqTCkrl2Z
KBhnSDFYtTNcmWcREAg6RebMxHdA1U/m4y+LhDBFfV31js+m+Yl0ymkyKqt9xoGRY3FPzXewjp8c
G5FEFuD94UIRSXKZ4en2SjxAfwhOxaBp0kU7NemEJ92XhERF6nN+hGE38sGzKN0xoRe3fd402rKT
Dau/qcUL5hBaxAFEyl5pQFuzohdJkZQ97tHTqgPcqQyeUP7X/ylifR28J6Z7qcekrpYmmq1LU3CW
QEdGIwsJNz+3SasGou9df/eyJB2EJpTdHCljdy4mDZQqoIODZxtrpyqR+uh5KK41yZQBrzpI8OKS
pK8+JZZCKlvb2t1wYUbXPmKI9XzDQNJ1X0lByP67Y01v0lyEJf2na4G+wV5hTxLKxGMFmb5Q2olZ
6KnkAvnyn15CiLox5/pumdIEr6bc20e/Ds0lvq6ZwlC4XLfIPfUgBZJ/Ee4jHh5ke8YVqkqmvW94
wF6w9taMstIXOpaRVAgfq9SGi5mdBa2SOq7qJ9/ei2TamwZMQSdhiz0Y3vDZq41Qwrq9ZaQu2TCd
/XiPI3lqHQzBXtGLHvfjz+mvBkkfq1EiI1nQB8e4eX+6hi/Nn+ZvGBD6vdedyfWrkwjZqbPMtor8
h4yw51KjxxtXgecgk/wJPUgFr0TCDmworpMb7qlpvg+I+vtQntvNq48WjBD0mXm7vwuYsKdwrXxQ
hAp1bllqb3HihKAmtS51x9hNnDt15G26Td+7nksrNQ72nxC/qKs2JAE3kvISdx1PXyD2m8JwBjUa
rfvpCdC3BO32DppyCwrtFqx/s+4FjOENqZiJ1Uvtmtl9/dwRX/vFjbdhdhS/oiby3daz01YeirG7
YSNp6VPT2vxdnPeucuRKpmaR+0VvhmR41v9sGJ1ra8LfrHJV9A0wlDUfeBlbCPB+O0cZq6DOtCJI
/32dD1eGw+yG2qJRnIHp1ckwFCnos7y8GMdWBgxO5NiGGKsAZ00fkckKKpi66/S3uHSew4r+c/PQ
ik6vPxcQvQG7lIconSUJP3kiCQrzKx5/QY8AwEUgIKe5V93XOOi6bvN4Mc4n0N9gotYU6q107Zf/
byRZchrR0pGGPkOPIr27g+qAx17zyyYY9D65bAF64aZ38KqCgBeuFTtHe1zohIuTx4oDU6qGaL05
xNAc6EkYuvuFNI5c5omaIiNTlbn0FZ2MKaIFObMXkj9WDW7Doj+b1Z6lMba7Ys6hPEc+VdhKctu6
W+0YhcgilM9qlgfMFgPL2CxagXCEGbSkzP1cqVbYE/uP3l2oMNOTDT05X5h2UgjiLmCp2A+pL/aH
dtE8cv50qvo0zyWI9ySWiU4spXcrogdCfUxby1ojb4yx1zBtlLbvsx8gjKVupyevcPgW8j4h2ITK
5/ueP4x7kOJEaktd+6L/tXpGqjMQDYb2FWxrAvtsZeQK5HgXT40B97L1kEE2Atcfvlyvl+6GoT74
vd2dNqqWxs0cqI2rZ5l6rmTMNQx9ejSxhuIZRLXh3+bN2jX4V7WYW6kFKVBGzSXdSCDnQhD0cLyk
STYfmGIbrAIxpRi3MOmwLXY4xEmgSWgWVe4ExYMsfaxh4//Ifv77Z5ZXnIy5AZeCO3hT09zwd/3a
p1gAMYnivlPgtm0yDPHTOY1Zn9lOy2GWTRu/MLsMm8J6otme13zQzNRK6Ki2XA64m5rrLGrqzI0C
eAtkqgKc3J4F/+6p/2LblIeg5/lzmPjzRCxH7WawbmeCgHmnQiKqvWFlGBYf9eotlur9W3tQVkS7
m7wjSLmfUnD2Z8viXi7zTiD7hb3H5yWNDQSNBXZlMIrcWRT4hS7phq/OMGIaFfNFTLQMwKR2XDz5
NZCdzVxPmMTmgMRt2H9YDplpvao7JDkhpWMD/NIBLKqkZQ6D8L80cWokSltbCbE11U70AowOwbX5
qRkf0nVc37QkoH+Rkpar9R7Vwx/VC2yyhat84iYmKowx25Azs10m8vPfNEaVlRXUqR2j1KUsfel5
VMLs/jUE2nHrGgfXCXXLA+Tt5TnM85tau+KTbv4MZjeat/aTNQZ4aewlOr/msSlURojtpekQ3feu
YP9LKhQwnRL/vnTUsHvO9IwXrT66oLT3QL3utbD52R064zr3pOz0R3xGz4RYBDUBCImH5Zydjnq2
VyX2Cb2Xr7SiVjj9bAlfGWKEWWm4O+MLfguRbJSdpiND24cH9ilZfs0sq6huQ/bzE+Yx/uwVJ5ur
BUmpbaX6m+ce8AxFeohCpbTySo+4a8WC9mUjpyVdRde7X3uHDJzNHisTdKi9MFMFFvG0Tieb7LzB
JxEfuYa0Juw3SdAAIjY+avjYidQIuMrOxgi+TE+Bc3mZiD+kByD2xKAy6YfgP2KelkA/jFYi9hpt
G2jiOq6dxh7rh+UgesOVfLJopcK2YasFGjGWpuRdkfJHJSbF3zxN8VvL9OABuS1y5il+SQRoPTFj
xWitEFj17b528LWtT+DU79pZZJF52cv7aXQvLbO5XtZSM2ShHPH3aDG3JHnwNkTpDdipcG5B2pvW
Rdauc+Y5pHhwZ3OhGjoTe1855pgNp+gxDW4FU/SV7U27PO6vNVpsRWMJVdQ6e4HLuR0uhjpvXjR1
oM+egghhRbIe6qYTPqsr7beTV5nGIPxPWTvZgFIZ9edSKA6omNcAbg5cgZjMyxL27tYPd6ZFK7dt
zfAKtEYppdN5IbKA7emMp8VjkD2SL90ZFTbkCfjG19QQQSeERZ3hImR4yN6PFYL+tZoYtbVizqKX
RAS909DxMYygEfVq67TgftRQ9QLpbFfHe4nDa0sHfy3rrgujufickf3xtKaqPcI741s7knf0Ze4a
szgoHavQTKyee8tIuOGIOv93/hyUeBZB27q8YJED7qKsiUpts5yEkbYMg0sN/yzc7vLY0aAgZ7b2
RZ1Gqr2RRAGWIZwcswTas2FK0ehDufA60TwJM33mVZ5z6f9Nd10v1EJ4gFIixxN7yo1QUEVR6s2H
cRL6v0PvKnvh+p9JJuaKyLHVVV691AbxKz6Zj3Pj8s1EZQUPxw0G3v5jGsujttYLUWHyGVhKcGpY
LNEU0ni8dIgk3mMUKNGZozVc4Kfwx2kV2+8oM9D2Bzs6V+VLGxFcKOrAJWqm0RrphDga/8e5dxRD
SdlEr0Dpivgmix3HZuynV9bajPJaCHDoUZJaN1XxkT0+C0sm8XbZVTf1z+7/1u5hLAChdPFs7n96
5EEUy2mLyziDr5oDB31BkUyTIRa1iG3gQRH9Da6670nQyBvtLyOLd2GPBwqNGe2BovDFqd3SdOKa
oEenUD4fkBs0lFNzOiLkHjEXy+fgn7WpoFxVbUVp4ih+wlzIwsN3Yt75YVPQeFrJd5cnkTd3aZBD
VQZl8VDg++4J7PcA2E/Ojnxt8SdoT1t0FAl4yFo9btbCENjWrtf53o/oS5z3l3Uz/noKaf9nt8i6
FX3EbV8CG9ij6AEGol/g19yLVFPoeHTsqjc470B6yyaY27BJub3Zwu8l6xy71z4BSLuRPqaXcgUG
GIhivF9vi2Naha+3/4aPRDpC2IqLWNGLbWUm96XJl1mepKadnOWX32yCiu+GypOY8dh1pgF3KifP
fNwweM175Aa9ELfETFvI1PssBzBQxJFajlSwJqeynNjrLmL3bBNjuX0gpt8kYdQqwmeuGK/+z3vX
n99JMIZl79WijhKt+mS0RKQw1SL+J8SXGaIEWzdcraIEyKFIXnzUPiaoEvOjQDwoyqRETOXWbCgu
MVWjE9vUB5rhNXWR4oPbAAC+FirZAq4UzQkyz/1ukFQ+75AYO7fmm0REf9/9xx+OzYlgMpmjvegC
nD8NQV4uDrQ+ov9nA0+UcvgO4p7KZVKb2zmgvN59W2XKuDH8VJ3Z91puKp7iD8y6ajATcdcxmMH6
y9XMatetx7nEpUqjE5tCsfWDDSZeC1Hj9fKu4jNN/oFx1VNWY7yEcU4uTzWEFy3TAykq0Io2aDfA
QSkgH/t2GB7viqohKVbQoh/lPttAaBXUC88LmmMwP7P02UUcPrQyZXPgqj92oJ/J40iSUARwZRny
W8IvW9ZizDkWENc+l3KF/KWawcJ9AaBW7O1hFCMJGvAAigchcrLE41eGeuAsOyWdIIg8KTGcZPtf
IUUUEJZn5i0dXpN/ytO9mOpRRz1wXmpYN8qasxXfCqlpmzAZ0Hd41R7BSqtliXEJh79Ht7DP2QbP
CrooEuDMSy3hRWPNBKdjzpvN1v32lWQf70asWQ+eudNU60N4M8EhCQqOlbNenUfHQL7GfpfkRQWi
mJEZxPO4wOgfD/nDSwLqpKzmYat/4rpcGDJb3fz/iFfKlsLd4JTYkMSumWOqgl0T+e9Uic+0bI2l
hP72VrrqxCHmW+E6fBxhWlRjnjSS4RrzNPI2/+UmD/74+mU7E8YvnWBgwVaKgAW2Sl1lkSS5bhyM
W4Sxg+3lWvr+wIlGbg/wl4IZaKvK2/u+sWAKWiem7mvvBvFUMQJDWN4Vq57hCyVWrXkswEzpkSED
m4lGxbRt5dzsShY4KwuRzMcLr/V2S7zKXkFByymsITv+5kBH5D0dUPfiLTYGuw8Wlff7bCtdSeby
YfR6ucQUEPplnZxfYDms53I8AvH2O5dNMcLmBcvERgdEmh3ilyjIQT6piBEGccIq1wf53dlzIO5c
nGoatoSl2GmYL+lo51/9evCs9+zcgioKmSHX9+Z7it6d826lGltXEOt7YLcl4DfiXCttJ7dpdbd2
D1fP8nKw8IEZcacN5jibX0HTNzjkYNYQhBAaoE9kRCltZXJSc/twSKGq8kmlDianairtddpsF+x0
VHoeweUl+ueTlyGwV9CpIbmCv9xJS3Miv5lapDK3/19WafdtR6aFSRE8p5IzUwmALjatTuW+c3ey
L+v1sObcMqzPr4V3cGCYZgiCAAYsFxSoUf/mKWjOim4F3G8xPWMuQESuKnt+DzaeS96aedP79XwI
yaUyZBqaQ3W+6qVdTd9B9TQS/3WmeI3AQesB4lijl2a/Yhw5haDWzXYf1p7WxS7WUNyRgk55VuMq
DlUSg3l29+zYEU7TDIBAAb5hPlRGc3FC2os1B64qKWn/6RN0FrPTVxTEwGUyS69WNe/NQNAh39xZ
VsURgSzLbyPINhaevDzhidTdTcmDjppHYI01K9IhyC02r4m5u/6CLCQCQedPRSDcjpG7aXyY3RUe
n9AO7tflPe0HG/+HRexAoUvBROJjDqY2oGemcmahTXE1vT3OAi7cVeBCRyVK2g0rWOzhAMid6CXK
RgtGZBRrpBBknINh/it+QVBHmaNhnzvp88ai3/QsKmP1n+otLzauPjzy/4VM3sTi7E5CzmABXg/s
6b3OCw/kPo/uIki9P1BsACSo4/lODxkJAJOj2PowGiSoKXjCuag7iIB5+OW0B+ViOJHaSHsJKeS1
+ayCackR+hMJewtdfK+CHwggLDkERXBOkdBMSwNGJ2+K8r45DvklGiZVg14qVvSZo8XpdcQSgj/a
W8GF7apgmvfW4QAqVqmiKUl42m2xhGjCN8Xs5A4DRHMKbbJITwj2ewTmMYZdCVlkcqekFyCMaTdU
LKl355z33c0FK8HSBWj8DpTHi5oo1uSUnb2D4yDIY4VAh8J03zX2saxjoZqxP3TJQ0aX0rG7VX3v
p7hp298ePIpv1Snv8fZwTKd4tkyD9PsyrzQ20mho5saM8VCtPRT329iJbj3UlucJogtP8JzkX3DC
7jL6HXRgyDTCtb00IqFlHyTXFYthUEvklQC2hVH2kouBq8aAct2VHwLx3+6XnH7oyzpGwvAxKPp5
Op3EYw5p0izKVOskuQntBStkyDbq8E/2/5fl8oGhszLO9NiZ+A0DZzOpMjq/21+55hO8LIZyIlcn
0f23YnobB2d3akC01MUNRu9PdDKhSIcpiu6CJMAJM2rRCPiHodKTfhCGn7/Ic6WpTKnoiY/Zvz5n
6nqLlQ/1QZEitmQtFRVzmaGiQ94nU8s1v5XznDEwHUCyadgzYl0hDTVM4s67nFLG3K+BsKbhnP/A
Ow4U51U8W7UZSl9vSU2NlW5lgvFblR0d0qFdqWFo99vt6irBMavYCphqc0roszCeAzNxWgRuvXFl
29wykr6rB2qaq3nhQ3oK75/WqNmgJ9+KgI4+fJTqGwnn3LCSt3gkqPEu4++2QETsbSehapy8CqSO
aYbcwNWi0FRXyiSdkHJB9oncZ8y2/XbR8YZKRqebF88CyGqanWxd8L1sZO+TUzjY9numURB/R1EZ
de/YfwvigNSqfmkTKV02VjTlFQn6oHCVRMN5zqAkFPG2liHD0b7zLgK2JATHfkO2ApUf8kJ67zNu
xkwbRf2z1HDIJG9TmQwBeCD7O8GCR0tzrpcsx/YpRWjQx6jYtyU9IZm1arIwsbcg00BqHd5/9NoQ
h9WAARImobu4URX2frVLdLfBJKO/FfbdmLUWmxk8SqQfD22aw6LCeDoScnZojDi88SFbjbWVxF3p
4NELUAZSNFodX8IvNVEOeMbqfWJtgcq8wJ/B1g+4t4jffVAqtqw0KkfIE+DrpQzKajga7/f43yqh
tpgub5HoYk75Mq1VPW37MS3egHkQ0hGofJ50pYhX7s9itoNhYtMjOJLLGC/1OZXBwC0qWTAIQOve
0NYmsM1KAXcdKLGUrEnHkijIMvq0CINbRhj88j031evIp4l8x50/Cm3HUKKKSQfEzUlA1OJQtIn9
RI+McCZLAO3vKzizteudY39RfI9rAO7pvcbvToErLXSxU7DLNB+b506ZwcFH2e0HSlNsyrf72sAJ
vNfuwnAWkeVCnlhpXZNsv0NlsQloKXW9ABv7BtZ/RyMreI4Z3n7pkj9+5HA96LczmER0jAIYm8oL
gcom0Ba5sTM0iT74UmOkcFSFyJ61/qdRfoGo7CjdvoFlqCzCC8NIrVSCGGoi8w+MNKRvMr1TfFow
odLscER7duOee+kPE8TNifCgHq59f/b0FiJqkRlHgSxLYEIYHgIn/3TrB/R5sXisQxv8djqwDK/i
0wIK9W2tGY8OhbMSedOjqYm+A/+aRa1Ao3aCG2bl4JcJdSNjxXXpKXiyci+BjsSZSft9Vs1EJlOD
Aiw5NzL0UEEvGXIzMJSJuqfABhL60cI5SiRJmpheuMoKfrIvN9FQwWbTGdia+CzMsft5g+a2U8hM
ZxLbg//9To4xcyhnN6bJW8UZnD+Xt/DS5MX9kBe+QI0QpaKjPgZiJM/l9DpYas7Z4weMbO+b/UTt
NOY8qCSq41goclQzaIoYCP2VgG7ki8tc9tqgD0zbkH1HC3+suhy5z+13uI/UjgGp45kCn8nLDa7t
Wr5RMetFe33udJigZCyi4+WWHyD0CbUNubHvql87uLjNkSwICqSUes5VfmMi+g89xSvS5JaJsmIr
UcPtVGgpYV2QQ9BHaZorAAUU/Bfc1qoTD+D21BD04undL7mF1pNbB/GsqgTsGfCIUaMzo/Fr2++E
CvLSFw/xoln4Gpf+CHZnt/a3LZry+V79/x4V75ZEdxwbZpcp3nk5q4tNoKxF3VLi5jO7nrroxJ8b
K0eeD6LydioM5Huf1ucz8ZZVY1EAQ3bKHhMnyFrVyw1QEhiig4/cQnr3GEHc5vrPPYPdPmyfbP3W
MVtCNaI70mAakr4r43+2p/llE7Im56uk6Gau9zriS3D0oeqIFYvN5YM/GBu4x67N0/WTKasdvDPD
4iDz6Rs6JniPPL2bcvGqiIrAeSOei+NFzMA53C0XBlnIUK+HPfIU127noQ/FUxjRE9RwBJQZ9UED
MUYAAwxkbObP9yGqgASNejtWFx7wHbmXbWXF9sdtmwMTmnJPIEZOWJ4wZAkDqeI7iPbg2mDunb8o
FTXip6DKGH+GNMK9XAulYFwTe3HwnUzwgEqcdvWva9+GV21TnTL1CarLbuP9MgDGCcSZPF7BhkMP
gHyQHGo3QD2ASKn64ToNmjbF4hdSsDJoiKzrR7h+OrZO1uH4IwY24suPbpA/Q1nPboLGEYGuLkyV
28PZTI6ZNPjGB1hUJG7zMvfqNpyjbncwSyBq9dOtq0WxeSG27so8cahpKDPuWmEIDtS7oL5mlXtw
FvpJHWFvg8I4pTjvo/Ch6rxl3BSHKUATPYH6hFXkF7qko6dDAQCNx8Mszbz5IboDAcTNWxirCpEU
Nps9u8q3r6EXsNJ3eGgnZ0Elp0tQiy9Zw2/rR785MsEusHfVJagDCjUYo8JaWaAhREXM2r4+KBvB
klTHHiYQt3KJV26yceZZ4NqWgm+RO5DInoPHOuQx3jzXbzhOT27ePTTu380/qmSndnU75nPI1Ms+
DHI1Ks1OeHZfE9z7iukzamN2J/H1HKmFDphKf0v3FScO/JlF2GIN26goIEObZS3uBhbIqgsd0OiG
3slgqApY4GbcglPMLR2oPOW4rDcTu3RJPvfwO5oIUAzNW0KdAQyxp+Vz4BkellEooPXiCuwvKpT7
ved/fJgYxNbcgLvj9o7eDlbKdl1dRjt8TFZHhvj0/1hL6I5mdgv2AyxYBhrrXkg77Kd/6Zv46bj/
CP9mfAfvUzjVRkJqcOQW5Y8pQ4t5VCbUYlhulxi4eFTaIEaFDa4bOLe/o5kRGUlwyTJv+N+FpVqQ
YDHLDOx7fvvABHQArcVSuvI8uHRGz3MD1Xnrsb8cregEpVNPbFxcf3LhdeGKNpT2D6XjiP08F6Xk
JdDTxmAJKQy3nhWZEwn//7zBJCV6Y+Fl558oChhRepz16lRX7A/TspSXuDM6kXWt39foUyOPsW9v
J99e/S3cX/zrRc9CoJ1xFg1sSvsjABv/QG/ht0OUerWDoqtWsyq6v1BeT6xzZ2isc6n569kRkQwA
SPIodCxooF1MbKGImZTamKxvKffMiqvEOPEFWs7LHBZI22GaJGTUNAFZU1gMfGAbaYyKNwg9AWTV
PnCAIPKNzrHnRvzdkDudsTBfIiRXCR1M5v0ffBxDKYg3TbADQBP+i8p6UWKiPnXQvPBXCXbyr/UL
Gcc+gVoZZDF7p8GTB2vKtAXkjgdY+MZoiOrYaSjLuHskt3DGgxgJytPzLJfLi5pEO3or0FCLocPV
dxJYD/2P88CUaNA6X7C3pa7Yc/S9E41EqkAH5220wZw57hh/5BJLzP8Mi5hTfNXhei9HwsKoNI7h
9ymQrIKAV0+UP8KRXxPHSdJ9MBQVUI4PdUIr2FUefMW5FJQNNEeqrMDptQYxT+3YpQWhOR09HZpw
k8EiK+4aH0ZIJAZ51llLR2b0aIo856ujE7tW9H0R3lV7KcUDpvEg95GELvTlfWYg0xmrgHoUtjL6
msxj/3f90Qq9xjOg5gZ4W84tLESGHgwLAAhRt4DYd661xBFpgsdhha8SO0QnoJVR3VncLu02LcpQ
djulzN/h+0pl2hbUZWfh71ULLffG0EID8bc1GUJvQxlYeUouf5V3K4nLsXfvYPgCDAPmD0XlDY3t
mu0LiolNRqt2QHtzHHKdg6XbRugiscTHfPXPvErU5ocT7wdqt0yV1gdrYv6Ap12GPAlYEmOMMeLP
MDECBZyz4xBbKbS04KO6OkqeGRD8CsOYt+nILtMzac0WksqQwP/6K4/IGARyKjdxSjHF3YOgsgY4
V/mx+2a0f1rzhXJyW6l9k11muGbfvtDxhht37GYcxSFtWcc6C1zP34cHlcrQeQP9+pil+uqcNe3D
6RYAP8Um/UiV7qwsoMzbe7CCQ8b3oEwmpkvvPbF9f/eSZ75/mwW+OdsXk5v4VeLcq/+fBI8XmNX7
oZemNHr1QJ260VtZ94FYgoldBdNIgdaswEKPl4oKc6VjFow9fixqubV/xdwe6VfpSccuYfCvnBfU
JY+F2K4H9IsrPk6IrRUrBRpLm3W+Q9ne1BLHkQxE81804tR63wybdMUqTuaRjwC9J9UuqCSSDCw/
Qmlt5/ZgiOvHX+lTcosRIgzN06/nrnb+agaPA1zYPzOjpPz8+yxm3d82SDDJ8T+YTmlkmimbqwPh
KRL/8Mu7oHcNUSGk1F1QDW/jRS1/A4NI8h4WCx+CyN6a5/Tytk433AgmO5a4uV8OjHa46TptqpHu
4Y4pzVk4bAAHhq+YptMz9cVl2x+KUnZs1bhp8qsPYxNtcY7uAj1TWY1wibI42RiJs89Be6Fyqbqs
CjdjUYzQ49uxAGyM6yiNQS3+NQU2jj/0si/4j6agvzvkSPC/NZ5KavVjNFExcLkJv+kspgBCGcE3
15H5hfU9J+n2MWLo7Bz9BHILY6HU0pc2r5Iye0alRLhkC7aCWbN8cBk6brgd+umqIZFpckClt9CI
AsrSLMoinrDuMFK7rE8mUwvwri9nroQclnfCgX4Et847rm9ofLq2Hllbk+CHlLywO6yMtNYJjQYH
zSmvBDG2cHwvrsyxk9T3dq74jbY+P5favQtH3AAR6LeFBFlgkh3IvBDBMN5aqO5USVZF+26du2uJ
CpfQkLMKmq63VTPHSvUobi8X6O/4MC8pwTSxqYZEbj1KRWAzxwZmWJQQnLc1GvqYzUBXggdEoRkk
rsybE+8N/fswktcXc3qreesbYwZxIXuHrZywch97WRYDlKftuN5mKF0QCOx1W0ftv89/VU1yMJUO
OE2wO+ewXj8TmS9kMGY00oOgB+ojktzhdquFsWv0oUBrY9K+ShSGN9DYNEDclxaZmGD/Qv9ESxCJ
RMRXTw0L1oYbXuMBIoQf0mQNoUaaH5Ybu/+IhD0CkjW8ZzBmPHNFzIzcJ85ugPHRImDpXhiqf5uW
x+J8ugMB+u6jEhUgdDCIpf4L2X0A0ts5Wuq8sOV+K64e6RhK7TNRIjllCus5Na21X6WclsFfmNZp
a3ti1A2A78rY8PnfaEe3z/wVLVDNxQmAWRP3D5N5lJVgqLaW3Gh5PqlnmzXBylALfU54lfvGJnNS
1SVXQe4E2EgpjBFW0bLpjhsTQN4CqGqSgtxKzrZU5D3isSdTgTES6tTbTRovWaBEmk5QKT4zrkSF
n1833nK7M0yJgFMXdyDwzo13/Z7SSlvosO26zQg072kbRLZjxBTeqKb/IiyNzHaWtTEcJsK1IYH2
kjXEppj/3tm5VeGe2f/DSJKNyVrX8oA8XImC7Muf2Gae8KZKREugDUfuuClKLpP+P01cVq/bJahE
GXlDuW5FB9ub6FZwYvIc9FIvSl30REmyLQ3d0HE4kCyxc2s6NfXYLGBqrZ5n1AWQJq49VDMT0oa7
+C+0YJIRbwUV4pmSZxkW1hNEMpqNpAH7fJcV0UD6uZFEZDhEwwYeWerqP6PO3acdxbBFsgJqXEIb
HAf9/iij7TBKeA/iI/BmqOlBYhjxBMDX2tQjBRDHGhkODVtMJfiw6bIr33gW3f6uKuoQQp4uW/j9
6fGzHMb+kQRW7+EzusFAXU1tc42VmBMtmgJ7lJgZdSb0uQ31s1HAcao2M3pHc9ctTue8aa6Hhph/
PuPAEcuGsihcLL2a+To/XPbEP2VcXL6z811JghUzIgbisNABoURw9uZWIN/EYJaQ+HVbKq3/DExy
q587Qj1+e1hEv7YuHMPI/C+bcpOwaEYx5Ze42Wz7TD84eII1vdWr9V+dIwtI4taHin/wzmuOngR/
QVQH8VGJcls1oQKDaz4t5MPhsBMqF+cVB6sfAJ/4KGEE5lHHEvTbaASk3bcFIM5U6sXEJSewI9LX
XEqQf35tX9E3xdZKQNMTwu6+sCiIaPQ9ryrDZ/UM6rO5XJq90N1Fkp7lnzjBvUlwYTyaKV7Lc3gH
9b7mDrKtn5Ewapc/k23PgQDDR66BuBt0OnekNFQooQl5+gHtWzs08h83eBJddxJW/PkSm4JJJpSY
U4y1okOTtmelTVHo8rYNJ7Wye604px1VUVdPC/VmO2NxG/iP0PVrEcho8CkQp4HQsbbrKuZE8OW9
rXFvngDdR+aPt3NLe7YTOTEhANa6B7XQP0YqgsJ/zCj+AMrRhb09WeUhl9RkzYI+y6eu8vrQTKyj
u/pQyvI1gvJRtoN2SMkXboaagO6BBUKSaQlqBAheBEJWKey8R7iemOr4L44yYBd194pH5ld+tslq
DUttJM45M+40bPH7Zf+3O+yIZSPxy5dGDaTIIznGCW8OX2GApTGMNxXbldQHPcIRnIbY933f5XSD
a7xHINN93a7YHblykUZoFieP5MEMNks8q+CKV1LtiSJcqk2wjPLXb5n89p0BDToQkUDZjcFTUjUm
zMSwhX4Y5M3+EKmhtG5HVMFNQj3ALTMvpJV0a0iJN/Fb/f8NqrjHVRiX9Pfeelx8Tphp45IwK8cr
HxZLPOBfdTYKPaAumRH15wvsqJEQYFZNJVAH82gvE9xyvZkwTzrxD9Mm53UEqNZIjWoaeYLeW5Nz
5I5i+A2kdgaTBYFThKalGdo8OQsAhxShOpbIvS+uMWHe4RaegRHBuoNe2FwC+b2QrXZ5Yj15qGjs
mSWUIc3j7S+hkDwbtcKM0ukAnUGA3B2YHyREPEW3e8I1sJ4vNdTyqJ1O520QxI2+LZe9TxG2jIUr
JI1XRaST0dZ0pYa5gFWiwg6gReiG5f92ps61eiefKgjj3N5aqnw7tydM27REogSSShp0hkJkltJJ
eLtwyz8zfIWuAD5PYwdAFcgK/Rx0KODF5Y8wjK7n/J49u86eW6GeCuYVl0xlz04YJOfofEsHGPWD
7lozydNs0jC4WdQJ/n+0JDgxRYXCo1fLdC+ETIs5VoNbh+syloIXUZ4ft/ySAM50dpGkbPVIAZmt
wEO7UQ9jQ2V0vhir5ajX8ZOvrg2jAVQ8v8Zk38zUNAluARoEKbtgho4LTrKmwhHVVgUfz25Ym2pS
zET9TA7WCgeZ2B3xFNRVooB+8vDWpcvI0ccxs9N3zWkpABqom6QVEsAi9Z8XGIOot21RaSeR1xH/
sJMY7K60yeBpeblDiWXXN4325aZyM4kvpz1tjcf46uovDPdzBSswcuFHCU3Avl0LFuTcCATkVq+W
sFI7gCgXQkbE36p8m4s1EOV0bUf2WzOasLYxR8Vm/PWpMV25enQJY4yIopoN6oYqN+hrI07L3m/B
o8ZkmINy9qExIaustyRkd/bSf4GWlRmbxIFe0vUPByopNTV+r/XEzQkD7o+Z5uB3sEwU95bDDlWZ
92CDE/ywjWbyUWiYgSQt6cQ7sd+Z823KjXFSfJXmCv2uHFkW6pte67x88QyUS7xD+YRHgiTQhYrH
M83BHlG31jZyZ4jWh2BnZMelZ8PZaLLhJSrrJhihb1nYEOd667QqfwgfB7pWDeExsHBGmmTlcqTI
n5fPsQMb7HR/iNA1vq/s7eA6Qe5L9gDOFLkiwp+BLBKomSdzg4m3Nc/gQlw6enaQ47DGKI4pyun/
q+DunOiTQmupzm/Xpus2VMdN8p8V6OZNesPGwJiT3aKhuFDAIXksGCGKT7i4yYNYhADvqmQ7mD8n
DzvCEpudhe3Qd5SakSm1qRfL3eh22O7j4If+KSN53rJZ/cGnnEjwZvCw78qdSz3082A6gO6SMQPQ
7ujc83ZT7iu0iBhbg2w6cnUYtQULzA5/D2D0EjG+FBTmAVuNnYiaa5mZdMRTM2oCjEYZLkHbdBom
z0SF1ey47IVz58QanrnLKvkQeWu1f4CaSLQyc8ngxvNbVSdDORncqQLyoji9epKDFfK+T/IkTy3w
NkNE5WwUhhiNwm3Zr58dWgHP1tagPkdKV0fJSeMCmbFZb6MsHQ6losmytXD+E++GnLoq2hnn4AJ3
atYOzZdN5TlEC4vQLHixGtgiE8j/rFIbB8b1U0xIz4PiH/bxvlE1fVnbv7Qfbu8RIFXkLRnYJZhg
tXCAlXp35RpIjpvlTYGaV3tOFQSq7wyV+IUDOoDcbhSF4LFJP+L58X0gwiaLVpzpSgpAjtnGRLxM
WyLV/bRccdJM9801uV2A52q5/PG3kRFc0Pc/sA2f1WUL/yni/eb+aBpUFwT5XTa3RIy0yCtr4CkE
Rraqoql5VJLzqh/ehJCb4KkbU0ZKQTENiQIJERtHaTVY6yT9QblUPB3O2VxCipVR2di04Jgd1aAR
DxaUJ9q8cPsVC0jLIdCgA+PQ74r8Atgb+m6+Fi9EZon3Drk5Jf/QEoKAOGIgudT7UQUocgPoE11x
b9IpeohoRxybEQE0nx6BH5tqM3PnLyY21Tqs0ZokKQ9Y+hRJhjD6mlCU9y9mAPGQaxBGCyFHXSVz
lwS3/Q8ELY18DgSKBKoabFID1NBdTm06GzblfZdOu3HcHL6F+qfdOLr5cjZNgtScmMLtHkCY94Hj
UIBk9Zv+oRxzdpqJc49aBNTdr0OmLnWPXv6jme+4G2m5/RfXOVln/TUmCfqy0IFI2mEh350HEch9
QOmdq1AolE3fxZD3wtD4LrX0VJdbz4QBHhBgrXDvvCINYQcY2PD5RRd/zPHgUesA1ylhM2uTlWxZ
G4VmAXcxNcMYlX8of2rKko7vVgJaPz5yLqRLQZuaj325PH2MQdkoAyEvJb/GX0I8nblYSCnYSh3x
w4Yg4+IiBPsFrICbKXCOKoOeLAgJpVmT/Gm7S2Je0TKhpX9bJgSiIeZC6FmxNkn01ddLvjU74bNd
OdBwh3jElp9/2Z/AUsllSTt+SjQW+wi6vogw0Io88cksSUMQA7yIByna6nge+tUnuPt7C9Aff5xG
3budNlaCQahubOyeb0SOM76X2m7mABAaGPTP20licmWl3MXIu6EDQxxxUAVny5oUPIXlgOX75NSD
f/+S6rNC/s/cfqlCr2eAvxg7FUGFuPmsmxKwsAKTDgMooCfl43C22wk4uddJdEw/C0ZCEfvXkrf0
Xwv2I51XFF/2TFHV2qimf3i9lfypIuv/oJwNhZsWwE4LguGyzzdhpMo6hdv8k18EzHICwNzgfydj
MT+4JCWIwKEiw5U5mXwOPJ4TDwGmxEkiPbvpU9Uvb3DMRCimZEaZb3S4+PrtkgWfRE2XFhApJTI/
20pPB0SDmo/fXg2F5uT/ghMTIiskzVQTL/VPny+BRgTHWO2T+CpNczmDg5vFGI5FHqblKIeqTcur
vCb+mU59Lyd9268GjE8A2yXs6i/wpp7LKoeK8ISD04lXdnTMWB7h7WNatfK+OA2B41V4EfhevyTE
ZcJZzeMGhHsIoCa1TDyX5wEfD05xyCIegY0GOSdpcYtilGqp/NQqDjjXUEAA/+4P4MiDWOzheZUG
nouCPopZASXHPJSgsa2HPtVa5nfkediJVSzYA8+ZzdNeerOx4k7F2rdMRIaQPKD03JtNMX75EcPM
in/JOmpBuJEvbf4B39gT76KkODT5pzyO9W44vQkjUQ12xSsfjLwxvnC87R5xNWqbspLWjEDYjreS
MLm2z6UjUUpQ6318mENGhpo/Nv/ZlFzTcubkoQD7mdH0d+UhCgFX/DAtPLgJY9QUlaicZoU9kKYg
qeTHlh6CxxyWgsb1CdDJWT1hPyt4aw4PI/ex5uAVeS64ixZkLQ42oDVOfIQHuXiu/DOlLlXtsi9W
kF82xk6UwCLPkXhGXPOJx8taGZZWvQs0eH5StNhMeE/V6Ggh4MQmEAu+Wp5nYZ9sG5Dx7oyDTmvW
s93fRHCRuNzE+6q3Qad6NR/fXOAIA1zv69VDvs9WNgfSkgBEqoXRqrOwGv+5947agQPLyAoo38oL
Yw/IotOCqq9+f+/K+43wacn2JJAhbE5IDcw+YhbuBEL7NIF6TPL0oHXA10XbMlWcwgspGUu48rRf
5xx2YNriLq3VxYfMIc0aLzzZ+70NPr2ZZH2TuH87kO1ymind6cO7sX+D+rinHQd01gUSUwgHBY5D
Gh6eR5SENPiZG3ugp5OTyWjKXYTbhU3QA4/1AUL9kcHG59DmnsxYMgIiWvS/R8J3RlJ+BtUzclfo
aFdXp7ix278sb8icwbZ0975NouB+U3U/zfIpFOosACHeIrwi52VE+qQ8a23aeL32HqCzpKfK+pwt
5yICNf9wtE8YqJ4Fxe2Kkgdy2zJhhI6iHyXyc+BYTHnDvhi+WbztiiSC4+P22G6tS6QU3Lj5Qe+o
cZGNvcNEpIj9mNUhuhhS3reuQyWoFxfLJq78PiBZfljyDTw+405pLHiXa3eTi3sNPYLTq7Gaix1H
H+QAR/TlRs1cIxJot/RtEv85boj14ajidIRYTfqFotBa+3kwkXNSasXv0CVGdHBCisA2WMz3pfj+
3t5GlEy/chbNnyfWoDjn6hMtNqxrRYdbB7wtTVelq2XafNJBxzXwf2r/8FNcUznCnIy25zvAiAOw
lY1WSsP+8UQ1W6uVtPaYDDL54oAOxXw20VS4IjLjbyTCb/mxKhatcaOUBxPvsWaLR+MVvnoBsvFa
uQ1XNSSAQzyzl9j+HeEAsTZF/kIBiWiCeEVGPfUEiPxtWCL1DuWMJaO/z4iellQ31OpBfvmJrPNf
XwKQMmsCjwNEuI0UsAVgH3p8w/Ry3XI75mwRWTPCi7SBSQEKC8jX5Nd3ns46IRC1GxhGmr4xKM41
7Re72f8ZwTIMRdf+8xDuk6VO8wN+0tIp+iiNcOLGj2b5ExynYc7XdcuLZuDpVmtmivvFy/Ivr/aX
WbZ8fZ2KcudupcGr8HvZBSHCSC5x35rTTbnv6SytXu3GOT9CW0VXhlLt2kpjoMCca07lDNPAAACz
txDX965kQGXWAcPzmqTPvUF6dva3fkCSwxKSWbS3kF6yfdDUk+/ss1Zly1T6aCBrlVsg2JzQqpG1
849uVx1SAXKj0a6jiWzoTqhMPL0gNRcizyofOv7xUpaIG7fHE1zYgSA2CcLTdYYNj5bYF3FhaHnH
u+clUPHj1CbKGO2Y9t94fxaGNMZF2cv7UhQTuNgPKJzzuvU416llEy1TH4j2nlsrdpMC22Byzjpd
cXwuiMV79Yal2kVis+ZBPytdGW6ToPPQB+YaPVlhDXNEmcm1gKsXYei3128R7i3fgIzTyWOOOAaT
VYCXm5MDYYuS+tA96Umu28L3IY9FasKQcBPMg2H5KiISU3HZeG9aZ4X2Vv6/D8/yHFALlASEBzGg
k7dQoSv0JDm6rAzd9pFsMm1/5a3gsaNypKLk1NESVtYUJyLR2yR1ln8+avEbMQtpojym44goHl+g
74S82wgnFykema60IjYPCQv339Bf+lxtLIiFQAwa7dvHZKvtQSe4mnnmltDYoyB6U2sXUbBU9XO2
rTmhzBJaWmQ4SnKoiJCPr7JCg1QyEhN7z/w+Ua2f2/Kw8Lz/AyXTbjAGgcVR3PfAE7MBUAONSFqk
JqrcrMhfkqI7143rTp73rN9ouduMihnP6C9DMa9ki3pUC854lssv6MZoTPv0FFkP3ngeRfZ0ILEs
Lm0hqJwhCFmnVJBfq6trDP+O+qVvQB6NDFxKqRO+vlBLH8xMUZSXKvscK8RCNyN/tZTcJ8gi0z2Y
eQIxDwKx57jzhil4cO5V4sn2nU0kWP8blrDHwew7C6TbBFzJJcLrN0dAHqr7a+DgSYeEQQwX21St
nsu1/NA3x41yzdPJWo9p2UzebK/iXe2GUf1rcme6qbmQSVR/zA/pzo4hTksNhko3KEVC1X15VcRR
d8TVOH/Mh1XUMeO5q1pcPq3oZljNg4TzeQMUrGbx+zUHWdYvD/dP05vXpawhmhtr0GSfd5XflxOZ
5R4Fo6XcQBv9mFTBWNC3O0UOuLto13CLI3hLj5/flNw0ZVaozoZdVxvwtScXvb5w+6F9wR+8OCMH
7WzPYItwFiTdbz+T2ki2yqumw8dWFu1phg5xZUb5EyH/ViB1ZasG7Rw+zZN/rwFGo3MmZl1xpTZs
vSA0r4GPpucLF5rgI8oLnHWu5psNvN3jkbG3gUgh3kvSjEsMXHcOHX+FyUS8TsqcQYt59pgK3Q3B
vFBobPZLZB5p+yWCVEm7I0MC9ovSlUYb75S0txBukRTe7+SlkhYJMAvP0UShrPkTmXfz/GwGIANa
BdqoprCRDyj2WZQQM3wPjvvIdrDmzi25QMYnLXB1ThYiusYBebfCCWCvzLQrck+m2nr9rw8Xh5fX
tJ1cNChbFJ77N+j4UGnmKaTl+lWhITeJFJSNXIPU6AlWX91ZuUmb1pIXdZaoqEBCzxmMcYb8vdV1
2pkTON2ijn42eGWtmqXGzOeEYywsJ/Iif2ZD55NzhzDC4+k6CmofBJcQe8DaJOoBe9d3KBlmpAnH
hZ5hkZO6AaNppEYp37jqUtEDoezhj2bAdpJkqLfFBGIjs2FUwta2KvExpKsNaKdnl3SJjarLxJ5R
VfvP99j1R4OoxzMy2V/9bqODbqbXXtOq7KfgXVw5XYYg+a+SpL06Aj0B5zJqdqM/rHfvOe34H/7O
dSpPfFkDKWMJdR2NpbrwZhKnS0WNX8PCIx0iIsjot/S1sCtxP+jZiH6GAwRRRmzO8ccdJA1vZ0/w
vJfep7aSHnF+vZtwb2OKcFuyqvo93gBCgUcyrbzBkOH13Kbo6ueeaL3/ScSLiOJpdhz7HcckdG9E
OiNYwstmmC3M0YfcyEp8YInlnVe0OREpm+5a0Y58GfokOOMYcXGdW78HSVQU2T8TkMuldx2StKzz
YiYvcKkD1bZMVBuWBPQQWxG0fm1dH6olRMMhLM8lC1PdItDIrvfOd0sfMKgo6ix3/XsXzuoRa0vS
fAYgqBeU+Ac78vs6zvZsQA/Bzftk6Of9hupAxl1MbxNanBDjL2IPhO86BBGlQQ31Fdcqj8AGY6It
1sm2UTrMHGD3xZdaUbE3pl2d/+MoZm8r1Ij2S106OqktDXScz/h7LJ9ebaRyM6T69g29k48EsApp
h1oiiyVWmvMseohXWO2K3HtV5yB0yUs2EKHeVkRpBJnRrpxhjF3NFzm78tc7VFWl8mZaMVYqsRtE
+WIOgC6vI8lUEvilfkCrfmFNqJ0asaKXYEHbnEEzSYl0wws+f1HPmPS00waC2viipeD4l3ouGC/W
w+NnmiC6rEudsxl/1mRMnSkbnNKq1ccIANrqYTm186jmlwIM+cIXOZ0108KNfBskKl75n7yjpmlQ
b6C6jvn0EzEpl4mOq5/8YiR7zkR22FmxlpsRyP9/ixmK0jKCu+w+xuKrgYFQ36Q70YCO7Va6Vncp
CLa+NjdG3i33Ysly8MW/1TnBUIkMC9dxpcpjTEbJP3+dz1Sp51Hu8PNCy7U3EeGYLKWY4ue7fzwy
DLMmQaBbvPny/oV0N1wvf2gSXpYlOicWeiP1P551wqdwiPK45jjrFpoihS1G41BDdy1CS2gCBCmx
9mb5U5RpVFt1piqCBZjktvi9rnZeLtEjbjQKs0pQ/1GlGdc33MeDkPpoO38z1Z2tCJMGWf5/R37J
kkOaogp5sFgMbMIG6WLIBxOQ4XWrQIHCrbmdkUaK8b1aHFcKUsVexnd0jhOvEqsKq2Is+Frbmxs9
jVLsxTrQbf/WZ2AZja9T1sxXIHgaJWOs1NGCRT+Z+cFeES24VsIVfbDNLDFqBiMBNwlYR4+vaJJg
XVXdqTkTWmfwlbryxP4Pd50yIkq9FWAlTPb+oeIAx6jJd5mecceEzaCStSyq8Kg2DOnucLCmbnae
/hffjWSyy8YyIdye2qU4sJ4BiTNUi+2Vvm196agaWzdgIRqtKkxRKv/78EFqJgRae0qMeYEv69WB
mFbbKB1L+j2yQrWbQ+I/pmupjluzBvjI3sfwpIRPrycBZt83LOtd1HJ+haLfSJUmBXXC3L8vOY8I
xfISDBAB1OR4VDx6YvV/uPIRPiMnvveIIC8+9j/jsIF0j6nHOIiba1Ld7Dcg7sy7Dknq4baXmkht
k+5rYS+APdL33k/bCWJYmw2PaOPT40kKHXIX8gUkOv7Lv5YzRAbqq4/yospTIBqki8RvGqcvYGuu
AGddUITUhYmh/u44Q7TPq5vA1kgVDoejAysKo8LXn5R09miKQeybXRxXr1X+vHMy3T9BghCpjcgX
CjmyDeDqAJpeJ/AWyTPXPPHdPWJ0GlInz1jIkCgiCWkjfAyN8WKyb3oGogzysEcC5SRwScGGFvXJ
y4n4aa2zhJCp3VbZraFhu/7bONqP68F3JVCaeccq9UTsQPYf5no1Lw9HYvpez1LKVvmEuF7ZufOk
rLkiEoEhpNGHS3y24cG0MWgSJn1t5QJXFTob4zDk+rv4FGTwDGhlPqmEZIBdkZlyvH7fx862LyKY
M7wcqBu1plMzHesXkfbiS1oHRZsQaazAN/xxFnTNIKHMluusHcS3CQyfHoNXUvk1gkg+KQQJYuKY
wGpfHwslbC9mX3GY/wF3eQgyxvWnXLyUirkLrDbbZSBnqcnjpspyONnsdLXCRB6Rw87WzvLu3W0p
f31CjGu7heIokxPYR4cod/WFDf+K0Rc4uTGWGFTUeT1AzVbcp7V2noNsWj13EZHR0rQSws9Clj8k
XzrXeiy7lVxJtJ0gTWO2ioqqdj1xtDAEoE5DfAeaam4sOdn5EUzLrU/uu+lU2GcsEEcYWJke/3i1
VDWm9duziNO/Grb1TZWxiBfOtUQZlQk+ojJRXRC4DuseF5gtk32eBK1WYRxHvzlx+6kFEb1gN7e/
WHcaooxcQsVqM1apQrt/X4EAJqsgbB+4E2RQpo9y2ezwDVm9JDNth1UcM3cxYz0eP/9NeE0nzlfR
Op8GKbl9lbI5DUqRW/zv6jdzCad/boahbDu2mn0dxB5l+n98Q/WqGXARRoByvp/3OJkJiDm6AH8z
Rx1JvvDhNXxRNCGnyI7Zx0ulLG0iEXIuNUPCXudmeUJw4sjU85Pch5HDwmP0ZjlmvE6QrtJSgmGh
7eMLDDwj6w9+yD3Ln7rw7zWCDoiFu098GA3IOPH2G0sgIscYZ8XyZdtv3T4RlXObObEaKF3JyEYm
eDj6x6/RhuFeWwqiQi9UiHtmW1z8TwbdGHvL+vHMXWkfj6YGeYzmDUMSAr959AiwnF9USJE7S4DT
+TccKO95HMJfVnPAz2FhwBn2CJQIQT2WqfG3F0hTDm9MZjT1UUoAHnU1Mauj1vca9b1Vmiyg/oP/
FfqdZzyE4dsu08pbmxnGoE1Q/36HVYO9t1kSFST4MQyb9o0WueJyAi4Bw8p9qh02ILeD9j+Rat9l
D8aDsKBBgcn6VI/GuVYX2jVaSr/rhFZe30NLw8M5sNstR9nSzeya3I4utaqOpJ+cyrTyKcube5h3
uyBdQgPolRv3ECFnJeVfzj7lkbbzHUzavDDiLZR4tdQqPPgv72jqQ2Q2RzN4JBxhPfeuZUhzAQlx
yq4WVh9It/5bQoY4Szn9ctE7BGA/loPVeuxwcWmiVSdJnozbQi/bRTI0+0YFU0M2Uu/Wi3Rz6VOj
ih1V81WsI8+IJefgeXOobvaRlqU1lJYguuyNcje5uuZDhPskNqMLzdhXEyrZpHfYFDdIsVRZGXFG
W+83wRe/6fIx7xFiHbKASkSLR1sRnu89m99b+g/2K11wWrbgA44PUtogBheJcN1TfNefJnaYvzin
3fO0c8/8LAC5i8PrGHYa7Lfvbb9gCBNBPgrDetxKmysXAY0mFBEstZJbjugGz74IgA3XrfnI8Oca
F8PvSsWYDAKQBN+7wbJwdJPqjk3UQ/VzqcBYIRocBsxKdoKozA2wAZCfQL/0bmGe8RB7QRfWiqpd
5PRcRmC0Uts2SyJhUHt37qH6KlW3YmRAsHa8L6u4BytV0E62DnqJUZNqVv3QNGgRb4QQttZ6n7jn
azKFX3WXbCCukmc+tOblKbLn1aZxlbHLvNs0BGkNXON4n9yIJ3BdVCaY6+cmf4AsUXEf3q+PxgOz
DlfimBFYk+4TtftrGPUv+HE9qR+5sVyaTlWvUqEWAYlnJjv0Qotj09upK+65uAzSAjQXsCGxXmlM
iuZKdK0FLYIFqRnaFSM/2H6BZ414pvL/UH8ZvlTEwL1ISGAcaIF+eNdVf7zs2gdsYwMq+tHp8G5h
2k9W2bWgxW0Fo71spfkYhIfnuZN2+2px00lfL7PvW2opW/o32VSygFovLm7+wQie02SXmWEbC1Dj
WvlTQLuiAq3DzG5dKbpTX08r99mk1Os+YWdTv/sfnwgbzyqag7FHq6d0dnTtjSAT23oqOn0FZzh8
1xgiKbWGU0GzGetbq3V9T9P36YXdD6KrPMDmhdCP2NjwULsBlnX04mLQC4H9qot06xdopcxxNlvu
hbBZF2hzqcgmU7IAGQAqfbtvaS4t2td7Csmt0KXyPUZKAo3Gmd8eWBJZOaif4n1J2ArkxUWT/mV7
kw8yA/O4cshaPwS5ChJtvdGf8UkhnmwfbnO+r95lgU91xk8o9VtR5dtEy4l7Uw0pAjNGr6b4bNTu
xRWZk63w1RmD4kCYdWnawMEhxzpLexXCjJ852jp0/tAkhhvltYI8Y40pzjLzl39wV8713pLkREGH
JcbO5CDrylGJigW8pm49tj+58lPLo1bvExqF7gvgsVC+sW13NkaFzZCEyZV8eXKCT5E7kLWzGEkO
k8HKyrHPgYxXwHGyBIE0rGkwP2sMyClhpubyFfIQjWhy+k+W+fq841cJteTckrTFKcf/HOOcbzAv
s/Z2gpcaV1t/UkJ4r9qim3BjXbBJQHOXzpCx/KyBlo0N0o7/rnyDspISTFWhxO1Unu/TWzaFt6Ug
vDsSQ+TPhmlH8tvPLXjXlLB/tMA/9u5xCITq64Zelp3HIqix26mOR+J6ugvkxXTraQEegQGePfF1
4BdX/ApZ2MKGdEiAGXEXcJypuKK0S6wgNVr7MPYjJqJFPQx9SnhqpLosOa8R4Dg4Sp2C2fO6qEOi
FXg3JIbhSvHirA2hgV8PF8TwrYyyXSGiLz0DY9M3xtKhL9ELzTDrWMAiclWF4NecgRw6NhUig2Ip
eUuKIqN3/C7Ow4YDeL13a6nGTyx8saqYCVY3z1uhsOttUewxvKR8xq2+9J3rXEqdXD0ugy3zc7iF
3SotA2F0fz/Cb0gQdYf++8MnTPDYFQvR/5WWz7kA1zQuK2icXM1AKoc6S+lI+SfFKGU/yuNXf8Ph
q1lw2WPaq9s988MvDql2meI/wDRkOSL7Us91Pml/XHy3/lM7n8pUsCVvhyxMsKC/M6FKq0IK82FU
VbPq969aahwjBnAKE5q/9q0MBEeDRV8PHZbTv9UpeS2/5WlUjjWC1UU8m3x5IYXDp5Y24LxwGb+d
C4aK8WM/AuVRanKnjxpJts8FTCBUWMIkXo6bOzkEtuPE5mnubZw44i8Xr6Fq8DO5jBHb/o/AWato
xC6zwqiAtqeAm2Q8NxAUcFej34Ls2UCShVIp/ybF0RjSe/2eaDfhmXAbXPurOFg3epDKHoHvRo0B
UUj0CbshQwZKONGG+9mTTug2jRLL+8vX0x7PLG2HzlvZALTnfWJhxd/xB0EJDjGcNHk2FrIDJxRH
ppDmBHtM0PzRiUZEq6vkGoBVSYVuDDL/2P7vzoxKhX7HS+zOLQB1/kqfLt6oRU4FrbMSd2oMUZ5Y
4bEJ8W8mHDAjTikKzcJ/vvNMHYSA9brPgqRENTULlDcxyJ2e/qKsm8EKLhyZ+/0GZKIFLnhmFrtF
5kUpVXJAk9y+xVeRWTGX0z+nhRuVNBFJWvVR7SoZRBzKO4wWWaMhS9eIj/jk0b/zTnLP9BmOR9uN
oNG8nhHDk1tUMYaqUmZ3I7uyYzotrT48S8+pZqCO+cUFbSkodTOrovsnEVajhM4U3nLgukXJaHa0
c9mBeND/oy1V/V7jm4888ig4hH9lAivEWLvGTbi6wUZQY0CoAvgE/VMM8VF9EDtt4kpT1kxVIcw0
7CQbE14gLhpzL0H9zsckGW92FC9oRXUHnZdOgrYZvO0JbMkkV8CQnxgGlK7IDjg6J/ubjd9O7UYS
pZODF5Koqjzg+t669ZEPiA14VYV2HOmMAFmabcyh+dOmY4JZ/Zab8li8QoUFLbJxETi4M36qozQF
c7/ZTBf86XDbmzRhZ6oQWGWGYt3/ol9iMbL8GIpS+9Wp2tMXloUmS02E5on/M0Jp4mP9a1QC8FKw
Ar64d7NbCj2Y9PCGjhKwGBx8xVmdKomxvVosfLDkU1/QBlLQ20Vc+iZrFJhSyeGM0YHZMGLwPM69
hJPWS6X10q3XhkFxay6j7OkXMZ22vFzXqXT6us+30P2bBg7pScJUo9mGImHjUXM5ZItGxcL2Jq08
pOpf+BUqRgodWaDQ7yDvbl+psmQnDo7chbdIsWUZ9hVXhMJXGm7WnmgvpB4y/UHJCRDdjBng1QIt
W/ZtAmiMDSgdeE0HzlYXJN+/rCqJKIQwTr/lHEdRK44Box/m8p/DHwUv4dkV6Fzhk714sHuspm4/
Zikb6kt19s0LWqweoay6gfcXxuWrkLi01QIyHe4RgTNWnrqh0bMQsujV6t+78wvVrcM5hqPqrPiw
HPDNXXYYdtMb2UN/EYH8SotdGFmLcMNM0F5mrAmvdZtF3wddDYca+xRhBLHTT7JgZdU4GhT++1vM
gmRlMRn4p4PKJMbrWbJUSKIDlV8ffTKIdcGK2qfzZJ8UWpQfE05a8udbRLkFd/6v1lcPphkguaIq
jlwzJC6nIjzVHoKbwHiNaunySWNfBXb+/f76hE68UXZw1HDAOWTFXChXGiLzNO6mVR/aVCzL99O/
Peiwii/uTIZQE84s3HY79bJTuxD21NIhAZkdGMOI/shFBIBYZ/aiRs48M3igde/nX6G7bi8Uhc2/
a4XDtHpuSA9GLsw/oL5rJ5JwjPe1bFZjTzDxbSsId3vIwE63MFbGO9Xu7BrrTOVo5ej1GB742dzc
oQml5LYP4BzSts5YGbGeRdZJE1pbK9YcqQjeCRJOGA1ZCQuIecJ70LOJOUqDBKdOIyI1lsZpwNDu
KBZcM1D3CCcDb2m7nhAu7jbr7YOs794DnnYu5EEJEy6Xv1DoHzVQU5P+IFVy1LirW3SfPzDKKEtJ
B5uhJDckPkNSnftBWqWfu1Wch/eRcuWGzQHlHv69tRNUHivWRmMn4MjuuulOBZmAyLwDSJG1tVsg
1Dojsf5pyAzUm+6d/csnbYjsWkS0qO5XGDwtxHdoyTkY2lDkQEWZnpesJdyPDA9ygSCaJ30jQgFG
lUk1e6Kmnp7jK+bYfc+975BJNWR0uXi6Hp/RZjOS/sx99359bWQpr6fn7cynN8eQus9HmxNb6uQz
R19l5GV7x4/OcCxA715D+aUWkbTBa/IkTDNm+GcZN7SZ1NFRguhz9KYT+8vSOu8NMTz+i/Jpe5vC
KpCm9GboBIV5jU+i4FVqPEqcOJZEkMNiZo8zIx7TCs+CiftThAGkmxraO6dcfoQELYYs0XrHF/NU
4dBiQ+0jZMAiVG7wdjrL1MEqCiBLoXoqSl4tvarp0LMEgKyuJCdyaaQjNy0D7d2wXH3IETVwPpl5
oZZkmY7i5sOAd5nIBzYELYYe4EQ8CHNR6PdN7fnCrU12CaJ8CjlWJo9zCMmwcF8GmglqZOJRZKCv
b5niNiy9BpexQ8u3PIpWOxWAkVb0aZe2qaR1SH2wNMoxkmv6ee6vp/e0hv2cvUFZwbCiouuCGEnG
UakohfDvz0wp7OMYgAU7+NR/9AyImv4LNX+rQhF2J/bVBAbu5l+s1T+fpOUeER/7IUXR3Qa5f3Hp
yRUJFyd3qMN6jNMfe2nU6Z98KIwg9aedV27it1d4uaX3S/97akYOOzIkiDFMlqgTNnVKyRP9XQOe
bdnySOny7tmu1FiygarPSNwaqgRuYpARP3cAQj4BDHoyjeb6wj2KmsuZisfsBlAguFQ7tQGgtXvd
K/30/Bq20AY5Y1+wL7Gae9erIZ/H8T09VeakrMMkoM8X9q6EpXIHpeUdobxofTlDQ03XbcbxFsMs
um4IB9/wx/Ol5dfGw/8yMlmE5v5qIWkM22Wl9CPHpnMTy0KBafQJLnUTRC1D2TrqRk+8/1EbZhux
c++snUk52LilyO2v3TmzrM3K+GcvGpnU9QhiyCdxoeDCrHG5sz2pzHPnaZwAVtWYTxrV3KYtoraA
+KXyHeS7drg4ZAbqGEYqeCzxvoMcOn5ldFJgRL6bxd0jeb0FDQ17nagKIGfq9uPCJuuCUicC/iB7
W9tqOpWHBu+kRRp9O2Y2EXBwosP3Uvvf2e00y99xXFOaxAlZAYI8HAK3bllxhInHj150osqrYJGF
isgUe8R91YRFSuIjX+JtjcPdiuDBXCP5pfvjCS7ch4glOa3y/HNd5a1reQvfUesioe0NurGlrFYy
yVSU8pzQGX+lzBDLW6ffcHU2R0h+EUW+XDJJmrIktpESLWPSREASzERQ9X6+ov6UtS+e+TGDamCe
RTQ/h0CN4A5OEl01lCYzesexivD+ydcQ0QV5zlSw/pKMqpwZKLXWBHvfF2GgMDYihPSNpIdXmMTx
ZwyKEXuFhY16726BPss1FD6DuDTmy4LrT62F0irsg+FYMV7chbmMHFHCDFZfhMpn9zVX1X0vwkrL
+t24R6xhdE/x8IiD9sp+4Mpq+2pl54R1y3rP5+BHyu71YaT3JzDqtTYCL1kCfJUqVPxZlZkONMdt
bdUaIk/85LSN6u96ffAfnB6SGolMyGWcsPO+F1wOuMWCuRqRyNVuS3DSskOWxbjSn2zx04Pjg490
oy94fKMC02WVLyhwomPx1ZJKU1ZT5J6c7yqdNiqDt0OFDODSwc3OpChC9uzubZ8w2qdAS4KoaRgV
40aQhFVWfxK6rpTdTAysaBdSvK3WLeMlDt0vXq54qHERmIFWJez5Mp1VOrRdKFRT0Ts7HtyCfnFV
kMro3GusAdLMKnGti77KAnOK313u6elwOnFyU5ISsrCoO904wo5JR4LUdGAEOOhmFqMmOonunGGR
KXoPNceoBtiqWQEztwdO/psBav1X400gjwATAXO0Gn8JTE4BPVhyxl9fHl4fRSlnppWWlQR+rtrr
5gBRNmzcj3fMr/Dlg32k3X1CDjoaUKbhkYnP3LrCF8+GSUiY/+886aer++JbQ28/KuiRZruS1Wzs
WWawFA65WanvndbpY3ljeZ+ZNTQ0rwI/Kk+y9c65wOIkTvyItyCC2/d6nXCVt2Z3KfaMpC/Cm78g
MrQdU/v5Ssv2FxzuOCfSjnuiF8uDc4SBqjK5/FAkyOsKriFaWuJA/o1uv0oddCfmIpp2ze5hlcl3
aNXcmltmhjS5pRIm/lm55EgGE8BaLNaaeSgIwKgfCBqwiMyyaxhyj9JGP//I7jJM53vw6nc8vDtZ
9iLpkYbjHfy7moQ+eCvsbsssPQlaIvZx8JPAnAbcriHwlKgzEJ4zjbBqS9ub61prmn4CmHzlxLt5
Z/UQqYfwTPvUwTsLZJhj6bwA2RJv3Q9c/ByMMOoxfIDLzV0lOZhe3An28XMxQM0ITs6Dgd7yyFyl
7N6ijxtR4TWgwVz45jd5enRFjbeRgr0VtP0usFpyjmI5PtdxKPIPo8de3D0Xcys32eCo3q1oA79a
ywwnyQWPiUZcqAFsaLwUplNNZy3U631EvbBXu0Qief+wOl77DfqRo1FcYAPrrV1L1Zc9SG309hkJ
bDhBQDclwddrRqTBHNDuFeYLMTYGo9mrl6ZELhDMkLZlY+mvjJfpj/cnw8hNqZxMFVsWH8G5pNVB
RfbwfWLEcHxm6kXLTGOyY1CgZXFyzix1C/IKPP+DT3IkOlwZ3zVhnSZsP4oN2RXkN0txEr5XRAET
w5NdVOBeJGniCuUGgSV8sgXUFvOSXuMsXWgg9bY/SG+R98OXjWN1Ot5be380JM56y1tOyINL1fPy
dhEd8c4Oc6A6Kr8J/fRJGEsEafUzni0K67HkueaQPNaDUpGFmB2IPCQNFkh/w+hDB59x+ITuMgmY
eeChgs9Qk14tvGlvfQLjHXij2AdW7CwzOuowDD1zH3sqn2lNSNb8VT15ArrEJu+vVNGwYANDrmrO
fUnvzC38PQub5p84hQq8d/cV8y/cD35Uoy2tGQemLraNbVmpP0lm/7rl5QTwaOKRHEpRU4hT7eq2
EQqbzJ7l/Mahz6Iz6oPMNvtA+H13B2LgKGSdWTgY24URxS44Tz2za++rEBZD7Fg8ozBbVSuWjNys
j48mEnVwRkQ/6mC/iZvUpt5SXc5Ps9UY5cZ9rbOA0f4ggGm3tvqfGe5wy/kQrxC36MFzu6Vqdy5O
w3FUD7cf1V9UmTsnnpN0FGs0mAzLYJg537CWjXYsDTjqldMVbRKO3rzT25Yrb9I+GL1cVWpDr81Z
qTSOM8h/aOgZdtD47/Tk9QP13XjSYOp9AzpWkim9UGwQG41QFmdL8H3cBHuzvwqDQLLMIFODcucq
1qig12Dj9bINgOW3IZlyFFkexHSeyKUWVWYm2Nj5pm0+XM8aViW7IQas5lezzt45dYbplx5t90gg
O915Wx58zVun/k9ob67fdZdpMJyuWv0Nw7xhogjEpv+f4vFxd6H5zrPx0kOWgPp5t1zf+xEjhAWt
Y3vcGF1CYOEHnUVB2LauiAJxoAiQ8MAWqRJPZVdwf9kqvqzizr07Hv80teOEJF061frfF4yxzOVT
f58GPAfpV8VjaO8c9d5JitAceyK4baAsuppABUffYL/WmK3sbibtPMLLUHCdj5UrLhRhnIy0LQGY
cNwoxQuoI40EFDz9vPufzqdKMNKyy8WFIq1kpkbVklA/lO4ZaYiZzBVNRazuyt+e3CJVPetqexWS
FpP7/4v3rill0fqvQie/o70J0wDzDE6LQfvNIoFQAX9ju4ufRR1RK5dvrdrxjyWf/4Jlbfq3H4BQ
+Nrl/+Lf5mF70pvJdI+hp6IAmZZEHxKczCxGeQDaxvLfaS8XAVdl9DaAINeXrvu/iaZ6Gwebc+Ti
RMMqvhIp+GXUq4faCbft4Gh9mXZDdfyWtCqmOsQXWELhnGE6IcfPBoMGBzJezadk88ECLrOrD4Uz
YJGEnickDWV3rw1HP4LWqsOIwYl3U64zXGdsKVDVCiG0woA23ccmnxUmjOkX7j8vba0HKowYuxXN
BOdZi9G6J5e12h2qMRcXreraYM1zQx2ILH9IQLNMLTYU2gjrUH3o4i2f408nBv/ryGm368qiuR70
jj2tkLp5j2HuYJ9tcFx8npQ/ZLwyW0AjOrl2y0HYCfrNjnNVq21T6qy6az6n4xf8zbPRIjqboEr0
TqrGxJa+coHoveotWWbmEINa9yrLOUkAnBmxPdwTpyW0ufH/9qMn9iKwknACfKIwIi51g7FZg9IE
15Y/kUYWh6aK1hTWgjizgMM6ZbXuX99nBK1C22rNgP6S3VEO9HOAvQn/mLtqlrxOeTQZGf3UqBGd
OeRvjDudEy1C/0y8If2rVxCvjlYaEzraERhwKp601fIHMa/IGaMgP7a2qdqaqVtdUhSj9kMFFfHD
d/y3UQaMkC2Be4fHJXZ055ihMEtEy7LAAXyunYdOl3h+/z10sgNZEvjnL0WipKizy6d8UhIfIGeq
DsI5UcufBcZVknEAVdu5YIHRP7DlFhO7Fn/sdl2mUSrodJr46CAfEAF/qBdFb4FhJSkR81tCGzEZ
4OTpxGuUlfJcYF+jd030GDnlelPyxQprwWhxLNoomxHlP8loUe+ie0uYevc4wYOdiBttI1UWfFIb
Myt8G5ob5Lf7QD7puCEYvB6Bjzks7D4IFE97swVacBtl0oLPQB7E/9mmzq9hJf5tbUC4jk9TjAnO
fevoi3PFCkc/PeUzK6Blo46UiGdgB/leeEG86yhm+DfYvz3hiSeG9EIqGib/6sDs2scX7KdDgpfO
kWK5VesCbZhZw3mDOSxIzdcUO8gVo1x2UR29XotNPAvz08haXQZ8W6fVHEKc2H+gYdftsz2pYl1B
swcTZAsIX2nr08BvBdR4uPhtOJu+igMLvPkr0PsGtO5CdjO8L++ElASGLAO4EwIAXapRmr6Upky/
584zEuuUV2XV855lxU684c2xIBFfrJy+ECIYOqbNjextVq3IkMwpZgYZuGHWV4OaPECS2eGcYcFM
TSfeTOkg33G/C1ezJ1eJjONctJHGhRBWKxp1Mx6C42xjvQrTlmYpRLSmbtcnydHevUwQ6OgnhVme
S7EX/cmF3etDF9yeg78SxxLqGmFu1jrpKqdrlYC+MrQ6y2lBf4yOfuSYyxFphQvd7P+F80atTIfh
mPMfo8+uR3Vbg438qzJkdW1vohl7/cN+BbfT/kPqHHT+z8zBic+zvKpm2dg78FnOthwuSWa49OG2
n9th36EgR1nSgMHYEVMlnqz6IszEbwy/HH0q9D6IblLdSCoRm1XlengarIVv32XWvrwRcwLgzltx
/PnOzimj9xcH+JZSAB2IgN9XBGR75Q5aOHTh848PH6vVMb3UvYu5bcycyRMle+advGauCm4KAU6n
4jJHqYZ9WJipOCAS9Gdc/t8+cZMjMHxD3Ot5pX+j5M+nA/uI50vg+Xai7qnqjBi9j/gVRXEJTRhq
mg4Unhanyp2i7fibDzGQw4B6QnmwIurA3fbV/seB+gulk75h/aimnZf29uHEBef2A9B50e8ZhkMZ
FSsnWrqbR4cBurjQ+wdKu8Ni3sC7ujFqZpprEEXrOhSLrOu4A+mByt+f667B8P9OXNSDLvGVP7fh
NnEaRw5+mcYxGg0r2dfOMDXKLJ9aCsYsQURsRJevnnarpkEAZZiuWJr2iV4VrPZ4UosNXcFv9iVT
u+zi+upqoA8HfIVeWoXyQ+92T2LZg3wEbBKmsTvPr81kljmxzr/vdBvbsKTyUZnI9/uUcfTM/jeC
6Uce0x3rag846hGWBYuSQ29IlRXPGV5IPjgNfxrIrCkSDUdW7f0gD81wyq/O6Pu63DLF7KoUbqlo
78xLxun+SspFBIZY3B+soe3YBltDyWszMUIdAHpzBJarRAFSAkbRwa/zEcHwqZW00/pAdWHdAra1
e/zaBX7lzPDcNImaQbJ7g3ii5USIVFfJTgkXd3rRLJqS05CAt8YNyQ4Tu6hJKm3puVe6Q8kkR8E0
Itvip3UoWbH5w28zCVw/V0fcDJ8R5lDYEG6+NIkNWhJGOIH1SBhpndDAEmGHOHWbr4h4YQ/cMIoM
r5JF+fj85OXMXI5+UxnzQTV2pghOpwXr+1bQsDttIigM4ibV8MIeKWzI64h5wn2pyW8q7FsnM1KD
MziPyguK80vQlIpzP2I7C3/TpyQC34kzRA2YcrysbJb86iln4DMW4LJYhllqkvrjTat9+YvlQtsq
Jsc0rcD1xd5naJLA1FMnkGQuulP/xlwOVDPpGE4DrMYPIZVtz8FUHa9BsJrSescrRseqE8BY9mQS
Pjoltz8k2qJKU17SxCZDcfB9NxeSPtcax6zg/vrBlkkzvEjA16wdIn9cfVWvDpTEqlkX5uKqYg9y
dP07XsEhM0WUY9vsbQXeawaoIvQcnK4qFQsQ1DMGRBLpCxhyoagv/qCZJcj5TBzzFPzw8wF0V8+q
780f6Um6pAkbIy6vwVXcgTfGv3pa+5qwNyCLD3Ah8H8K09BJ3oQfu5SpjZKxr889MXnw5LhSlagw
0dCNnf4AS1oDzWbNhp7k/KcjpPIwMXYP2/hNjSO0y46oOJFgGHdJFT6J86k0fXn3Ookzn9Xp404i
qdg+WzvG13afScUBZpQKxB+fPqLyL+MI5Ml4g57BZQHi9r1M1rsMpMxwUlveac+1LrQS/m6FXl5b
57SQDRSq6ZE+MkFcrS/ixv9K8whHywtQlvC9tbjtggHc08VrcE2e3M1QTZeEu+oWnVUywOEHe9nn
zNqqKvBB8PoM9eB5YHtbrpQ1hvjQrGQfK+quK6ysZjha23IFLUJx6acJYaksVd8+snOvLpEvo6jB
Kll6D1GB/tq8gGLU1snjLqLSOSd9dApYcN3eyi7w+JhV2uDxIKmQ/cho4Udhamm5KMHD3MAIF5Ov
zdBnp9BaMzoDEY2igACc20YrOC4ftRa12ZOHL0XS6Z+ifEej+nqUspP1fu2l2vvAfv7PLAgl6DNk
P6mO5vN6mon5XapPVv1hCcE0xHEjXyI01gs16XJA/2viJRumGkYda2TwVBWK5x7HkWpTPAni4uhd
UbeX3IqYMyyvXAJVWnR5+0FKbx+fg7yWIIo1mcIj06ZrWJpGAfjlDnsOIw/OVp0E4fAypZn+ygui
g8H14XfZoWbQ1icclqQgny+s01T0W3gKvrhRHqhRu4Ir7uUyUgaQWmkoR8nq5SQFhVEpgtP6pl0u
uc2BEZWeKv2l0zs+5ALsEl+8O54a3k++N8zLaby0c262YRBV5j0j2xdJlKvdv2NBULdWAOFWG6Rk
M8OA7odmN+lXJLw0jmTrVsZd7WWmttKy4N6kEJRPD4wpIPXrXqxAc7En2Mqn4ZcapVMc9wNuzrII
7VY6To7A7evmx4HT2fDt+qfZmpQQQ/Nr+cBtMaGoB65OHG9PU8+1wxiogdpF5YJKrKICdhuhoFLC
3c3lzgSHU6erR5NTN7aRHuZFalDoBmswUK6iWmyk0zr9IQdpuGS/F2ZilHBMDrZ6x+q2k9/OOVOw
0eTL+6ioBUja+fe+zNpBhONWvQW+ZoFkEhyZByjLA4fyXoZofMqJw0WltZfJrglIl3wbCqJkKTzo
hjJFHa1yLe4CB8nm7dkgKcXTLrDiIlY3JrmGVrIjv1IBsuxCvKPsWhMrvCjl9umPV5KN2oKKwbTE
Cy7OYBAaoy3VTgU/wJOOe5Z4h0dyMnmLlw4joTX4j6VETY1d9arKgIAPwTkoZtRetqIS4PquiWsd
plrHl0vY4dQ4DxufF89a36FofmjfdwOjwvJDBElQwREjm5gxTL4R2OxVB9zbPJxc26sydeSyHpUo
iNZPqPhfjp+7yznWOLkBSqhjC9l5fXKsTaPPpjbI/Z3xC8LSW4N9MZxPzV5bypOgJ5ETyttAAYCV
kf6n5ZeEVz+ZQDj13FxcW/wS1O+VaZGWtdVlH/LYfrLMwPwXQc3+Nrmi947Mqrf08cblqx5VPHtf
7hsYd3GlT8NaRqnl5FIQAdBi/l3YbGrGIbGp8GK0oPNUQQFhAosQzSqJGZcLPOe6kinfKdtfDCJe
uX5uJkWvHfBq1KWTph5QULFVg2b30HOdbgWm2cxPvphPkssSbxWFGgz/3wrf3fysvChOmbl1HnE9
T+Sz3njz1gfx9N2wpYEEALNEbB1qeIPbZzJyoT2mNgADqRo5aLpxvp8OaiUa3vr0vltCecy44P3/
XzrodB7IqfwnYXNt+bwaqQ6EuQqE6cWVtbVchxsFjPtobf7MXCQ1tq4mwEB5NzhNPN9qSUCHLzI2
/r02uPx+hns9sBJV92URNdZQRMeZFG5OM+bnCmDqp2ALywVNJ6Bfa7YjdE96Y9lmwHB+WBGcggBs
U+NqhCNm9adwrVO1CdpYk7NDQZdl1nkLGVT/owJwRFI42K0CJJ0UWRarP5HY81GMGT7MSjddEpDm
ZzIJ2Rv6sasj1Pj7r3RxlaZ89/JlZBBMSumqbU5eeR8uNuehsZGKtNT/4Kf9BzMBpUvaGLBejjJQ
q4Mtdgos8vIeoJxkuGQYUhSjLV61MSFENv3Ek9FDFQDJl2Cv5swL9GIJi7mJ0E8PyYpHWb8sg8YL
FjlLEZHuE4oohzxTdFsPRa1kXLOLhA2SjQGvRMNpgjd39m3bhMM+an5w9GNYh2djwKtEyN5NWZWz
uV82LAbwvO6Djx7fRNxJnUAP+53KyMNaPBhPYbA3/kXjAnkoIBD48m5zni8earIo8d4Mg0XxjA2K
V7ssDbHXLMbONOJSiUtWGkaWXz4VuuFq6H7+CeeMeucplhpRx0u27bbdFXeyZz3CFooWWl5vHnxw
biBxcj98QSqbiY9roHhQGfWK3dSTsXU27ZNG9H6nySxSZxTcLI/DHs+KuxaoP8lCC8uzL5TyTyW2
0dZpnjGthauSQpZrBhoGmWDYOYCxLto1syQO6sNDjpvenyb718HTfoRsNSnbH6yvbGD6x0ZC77aI
vfCRv/eqvBQAu8GIxDmaANZYfRSmJuIWWGJapAIZeUGfUNKJP4itPw2hLEKQNUf36QtK0jNARDIv
mGgx+CcqOH6hN7rDRhuRA0S5YTppDfDNdydrpWr8shwz8ikSDms40xJHKb+ypewYXTZz3NCQn7nQ
GXOvmmnjOgUm5LIavUAWJKqaNo4NAAmlOO3v2897CD3M9OqPMFAeFrDPANBJgbrubLw0rIOXO/G4
rIh7OzR1w0pKe5kCKMmM2/navWPqFfN2uoQEE2XkTqLDDqgAFUj9QXIhjgn2nPCGuwKHfgyMLfhZ
RaatILk/ryUq39w8NZuWDekjFNpwRrntrGxo1lxEteSu4E7Ge9KtJaazTrAbcppgPhKkWrByAaAr
fRBPj3vgXji8jp49yLDg4uX/HFplwhKAf+G7rWJoEYbS4T+6b+YgS90JcY81oXYCezuqwgxKC8Ir
kSgl+rVLerRdsjuNIlP5M6aGcDVtnCGBUQnWCtVhtL6rOehhZV9Vk77R+vY9xiFnfDE2GEptAENT
Nh14GtDY6cwfTeq2PyKQDHRmh6/wz3dWubx6B8ja784hWKzytlJvnHVAEfrX5KjxW1iXbKp6YIR6
XVUzJmNXhLyYW34J7YR/t844naUJaCUMkz1KVYaaX1aoOynx8Q3j9Odn+n3Mp+TYhmNDkAp26YTQ
x0Htnfx+ESd50KivQ0cjchm5FgrzXTetJyCqk++5uYOouU/RBmqUzvskWCbRAXnqJ4LNUCpFcR/5
aScRW1WhVKKjxQ2IwRfdLZp+i4Q4if0MAdv2brtrUyObSGB8kFqmYOKGaCSggRmPA3xgrjPR+QO+
1N92XigfIeKfhsYxE17Oj11mKW/WvNifKZy+X6rAoNhHAiLkksI1UCNc6Wo7/Ant+hthNgyTiOSw
n5VpGBZAleMJ9Eqg515KPL5twSgBGUvzliUwh9dSYoX65FS8VBPn6k8w9qSlEj3OIhf9ixlTC9zz
Jjlo1gCTsKuNhIciQCuSJnctqkxDpV0wYN4nruv39gVJtWDzO215m+tBHcyi5eSUzxTKri2CmUTg
on8KN2/9JwH1V0zwM2r1Oe+a/wXVtGRhCdbjFzFhMay5EGkHtMhe7HpFTmYWcZrfNzqMTJe21hpZ
S4ySCrCMRnBcN76eZHxPfPpBhNf07b0DTPJiKXRKVYJEByJflQ4c5R1ObCqePxErrZA3WiGaEZwF
vJHUi9tnGtdeqwNrMaTvZVUz4V2gdVn1LM8REt1H+ZlJhf2it3NlZc7LQ5YfAAUFfpdStT1Tjv48
RNOceyLPHIQQjXyp1HsmFvGmv/UvCqtAq8DgYeTiOLUjCTu/j5cbTTe4tyQGHOaYDvqeZM8cWOeV
btOMi/oJ6l3FzGoraA2PFkUtfmab64/6MZvRo15zJMuNTtIvBTNZzgsQLl3U/CqAgukzdig1N99a
y6VpkhsgF22+TOLPpVrsS9d01fz9E2njaajXC9gHhCK5gmG3S5RZPl1vBL6G3qiTuCuMwuTx/1Q4
DFT97cmlNTb8Svgm2Z4cgWNvT8HIVQKp07UNNN9neHRlZexA7EpgZRjR+xJD125imP86yGKhSQ7Z
fw3u8rz4Nu5HaLdRlFIwziY1B0zWxi3AGc/RWwgjchGY5caYgzfTnBqQ+FNJFV8RuFkV1X6BfuTy
mJ7ZvcJ9ai6ud6TBuKDxaKAsM61z0oCNqPGeUl/XG5PfSXQz9hsXZfeWJMBGUYlFME+fpzR3LudI
yHISN7mvMJtaJ1+LnfdfmlmpP2eR0BXRX4wfDpnVzAlh4cEx5+C+VzCol8EXnWI2Es995Zw8MjXS
ipeMtozO1Y+zsd032wR1YFjWnY6YQgxSBtSR3wPhSyNpuDR45IjlRSekrwEoMMB8AyyXe8UfFxm3
kIo1a1IWHo4D/BJSLZhwQt0vWVz6VGM5dvnngp+ROGvFYJ7oHjT8HE8qY5QHh0IzvBgu86PGOU83
MV1PDAQSfLq6QgUFm/DRQFee8Ms8v49x+nYh+zA94LfYW2fXw29KNFIqSEjcOQpksF446gTJddjI
1NCd151DBIkX6ZqZE2kEP6EckYSU1Lb8AXHj+H68KlvPiRxGs8Y+3FUWGAkvRfxl4dmO7/UuO8n1
ONjAEpLWcIr0s8xSnu44X8+a8IrJT0pSUf2hmkXg1vzF9s86wjuaPlQRAL23mGfSe9KXQxf6ifO/
89XS8Vw0J+pwdrnwKlpq9LTPejmSoj5ZCU/6SLr1WJCsReW/na32l7wiz7VEA8RmIscbR8NQBc6Q
qsK8G3ia6TbpMuIIKFpyLMP39lKFGqYpuYv4ZO/tPbFjq4FRrY+R+Quv8kvH3AlXD6wT09z4pnJV
pMRQJnkSPfGhDYSzdc63wP39K5HtFfdH6uysCYXgPy2RCeRgv4esOdVfA8a4rDpy6b3wCzRwaRt4
wfphy5vUeAnAuDtyahbEL3bs6K972OfpazdPC3lIhqQ5qw7EjSjf6xn7hmypcQPHQafxVEd3icxr
WNNmtKjHL0DyKzoOnsIt1e4+YtpVAArqkqpZhBKMzi77ML7koGn2PWvTcwzjirSsyl4Awj6G3BO8
SlZ8R+wQK7IGvysvagOKWRbbFmNApV3pEUJNXizrK3QZY4mgR/msROduq8Fmtn4pkKx7+p/sZ6Yw
RDbdeuBsngPRuGKBuCLapwsMj5RPP73FxRLmPV+6APEZuS6j/xhECymN6PQA3JFrWNaCdsjEoLTD
qGyfqi1VUoOY8MlW4aBeXLjpOEkHpWKZiC9JJRHGQucDVN2qZcN3vRfi3nL3r3Bf8x7Mb8RqNxId
gLVjLn3UTaXKiLvNC2lKd9uLQRBGomhFv1rzVo+LIkaKdFsDM4tXvLRM7SkpDti8asvuw2Xr3NWa
aY6J5fmtCVgq2NCCUHZ+Q+2uG0EoEYn41miR6gxNkkHBsLVMIRHDF2qIuV76Ban5E+V7LUjZlhv1
UZZtQhbl0Vy+zA/SYdjA1RU6EJ1xnmRQS+ek47/G+yPCJI6tRGA5GfL6LHuUbyzzWhy5Fk1r73df
IDuOMxQYmEVj9QHoxmhbAmoBCjQfgowIs+421IzldmzqmTx8k0d7n29pXdu8QeH1SK2+Aytx3EUU
a/kLat2YbZBo78i9OUX/CVDFMVrDroxrqFwuovkGXPBA48ZpcxXrEvfiRGWBC+SGh7qlsA/gDGbp
0mAVJNmV9TIZjPhNj/QERawxGWX3CM5u8+rMaq41U5wBgG7ZXoD8zOxOoLJdhHQ69AR501V45e6q
1rJBokGNKicDakNLITHqdzmC0He2JulclPqe6MGTDpWBs2ia/5LM0yW1qR6LlKriFjl11dZYOGWv
He2yBInGoSMYAZ/o8KaT3ceWaxjWivWtScHiGHGdMhIFokN0vL1LJC0gB4f5+5g4nLwaFNlkWNpQ
esmGJR5NXNjxiJn3khvgyBcIWV7B6D8qs/7eDBx9m6NrlyyqHdk0a2iQ2CIW0M9AmWgTGbFk1yDM
QWePaaY8AD9kQphk4XKL6NbGRiLxs7ADu5qPp5mEcIPMfCRDiCIXMfF3Uqt+JUs1DdwzO6JI6M8Z
2EpiBJe4wBmlHwEEolHzHZbJujNCtGeVAvc8Cr2dGD6fOcuk7V3cMOBArgg/Q4XpxUOUI94rYPEb
pCldZnjkwTYr+ar8gPe+TlbsYWac03Dkvi4Kh8wPzStoAvbj1zxKijMyKVhCMhmZoBMgSQFmhFhx
Ewz+E/9cGPSpLXUJhP9uwxKBwIwxnwbzqxNejW3CPcrlgt3dBUILxBa9D3MVSCH8S61m38PksNbD
uhLPU8o6ZBGt+sJN0RkkdBQPXdxZVtqZuNklE5ttzewnaC/LDoBh7TJ7Hcvx9jL6Sr67lMGYxYdD
gLV+XW86VY/xwyM1IJgdAVZejwWfUiKPfMUDpXskRPb5xKWk+R/3o3oeuU8PUvrXOdZqnoSK2caw
0NgtPCbG3HOb3FfNVGXjMWGfKVnLY/mpJIMT6WF9siY7RNbJDPgLfh0odi6hviTGC+jcoGVsZa9G
LN6yzjNNijlhqTTUC61ZirYBNFCyl2FjgRP0Opi8BU1GXYcMfUPW3mcHRIkYWPQB8NyPUOnDZS/e
SAolBXH868gPKmrV69a/AxIIwtsaYHze+M3L3DtjFtRzElsgVm2iMFGO9oSMSk0wDzKhRLhgJS5A
81gjRVPIVbmANe8CVe7vh1OB8Mjacg4QuuIWDRHHNOKRTHayQE+TNYWXX21F1GN0oEww5NoKQxMa
baU3Q5BfW+8/R0bpqgyI47+tP6HaoI3QvGRIW/MwVqK+Wr2yZl7EAGJwrCN2XIKCuv9maHiRFxgL
Eb9iayzq4TPj40swEguxvSDL05LuSj7Xpubk05x+Avk3oSkdXl5o3JDHqpgFJGZKo9oIIc+yc9PT
99UTDOlIcUzYrrhv7qKPiKRUb+mKVmaZ300h6uqD6B5nqFWcOlgI2mo0aPa7u8yCXlVq0E4TWdiH
h1aiSCZwLXbokYkBefEJM5fsjtc7E7H5ohuPrIg6y3UZ6CXWq6hC440VcrBeSJc5rOlyzINU5y0s
WE3hu5FGTFWr4SMJK7ttWfJxL7hsLrGDc4BoEK+H1BHza9Cf3swg49n3TrueolCqUkPvqm+m+qol
lrQoDHBhOHZFxRghs5jRciXEScqmeayvegB3Skg7rJy+rHLM8BrX556DHpd2LUYBARO8+EdG+SSN
AC5Moe/HPXokw1YCbh6A21WAej+eFGY8qWKYFeywVeVpYVIzSTOY4I1jWqbUvYAWLdY4OHnx339M
R6swuH/nADwTaudbcaHY2T7dEz0RbSYdTXO5YZ3DcuFGBR/6b1/vhjIdM1Y4RxQ+QC1flhJ609Yw
Hev3/X97NykO/irQEilmyzlKS1D3lCs8ejEEPHuU7ruUtamjGudFCK8AlDx7bsTJSv4SKRG3HZ5f
kapx90EasNvNJkma4ILqdFnyGo2nbQ9LsFhHl1qZB7cRv8vAJQYwkE332Buk5u3vR+l/AcbuobtY
ycvTlm5R7yl7sUhJCYbHswHQs6eKME+/ClOXdYZ393bJcDCvG/sywUnTfgAI19BrFGqSXvaNyRq1
ZLTUe06A8AIsEp2Ygm5b4SHH71MbGcYG5iGXYVmt7/ZkiEC2MS3Lgm+noV0quRW6yaa+qS+ZkwAu
TJgcyZPoEEmuLEsaL3SL01lh3svMBp4P2nS3ymZ9hcbB5tofGdTj63iAFOs+t1QB4n6i9+6Jn23G
DDKN+40V9mVhqRfQF/BTy60KpC8ODBfisezl2sG/PIFY8B0TepA4sXRBUTtf6rGJk9ifv9Ae1qpL
3+G/wKpxW3ACJEvtpOvH7EGrH4jqrP1UKx4cAKJjxdU2XLyorjsmlxMOJJqU0j6k0NPtYhhSFT+N
twULqPbPj8sdzQfwZKweFL68FnoKjOxnOtS3zxy/9YmcKP1RuW3yq5kdQWfSafUMLLCHIIFBOUCP
KSuEEyaUFNYp2Ug4zPKxOOLczYrFmMeIqnOMs4QC2cXt4vZWTY8t0o4JNF/IY8zCU0F3ns5GKnz1
EDlldQNq9DJuCr9ZdDd+wL982tBeE2hypb4UkSYZBjpDgFkNiZ+2hZ9DBX3xyJ9Z3HKz+CrbSskO
lqYKPUSSQlQ687Bz7Pep4JBcj8mJpXVfjUD3RQZReUMP/MAJVQRGrRlSOf5Y1XQmsTCImCUT8xt3
x9s1lRFvHGF4dag5GIp8RqW5oMu7SFqVkmaASsxQtTnOt8jusX0VrcshJTbqwRGBhC5W0TzLH2mV
ZBxCr5Z3j9quatCrufJX8jSHjgnIf+xhZsaek22IQXnNs9AJZGgn2dL1nfegTgDvdOVF4SAwSsfR
u0zqoWx4PKUuqRgfv1ICnlL4hlfTqTBT43wrgIiGVoOIW3bMbedhj2fMr5fpvqt/biTFfvcXiG8o
6vpncJ5dCD/z9owm8Ld/95MScPz3CWtkNed5vmFahpbdmM/k1nqkZ/mlacqUhrJ3zKWPpWrP6Vg4
5PbhzOMd2XG14RUv6HkLqPKDu28zVFe1t4bODgKM0IUuhHCMmeyOdxQNWlvgLESzacTb0j38sDUI
0PB08EsautHzT7Ou1GM7aDUKVv6ssKyPnL7t9NlLVdCiabFwkYorgn+3aEP6pFeJ865e5sz9K3gI
VY6RGiMEGp8Wu2WNO2ett8RFbgEhNWjOFupSgcu4vJfKxlWTD1jFOoNUJ5IF1Kyo+TrD5pfUIPOp
wmdnDHBN34FjQmB8aC1jpdGg6RCxtUzObezqICoegB+eRK6xsEgYjRtJL8F9NaylKFAzsUNesRiw
MIsZc1TCTeSk0Jgy81qreQC5qxhThG7Ne0fBAQxZO/r3lcH792n3z4K0ZHtKb0fVid4Ngwpol2lp
ww85xYj7p/5uCIFldMqo+xD45q41wYoKH48d14/zQn8+pmnN95dmOqPgsm3B5lbL7253631Mqttv
TqNIwvssKzkqT84O9EJjDwPj3RuU92d9a7HgztsKTWoiFpyZLRtZ6HHLrC9x7dsU04DdPufOLX1W
97SIoiGbVPvq172B6eyo8z4hsM8aai0IIL3DELc3nIOX7nP7VXr8GskzRoCLlIedkCnWo48jJLip
o06h3zbCWyLdgTMnrcuHLyT5X3dTIvCMPIWJGLanFGsrxyaKryp9B2ckrFV8zvrubtqjOjTQ/Uf3
T7YAAbbdRejhtSlVUBRy45rsprIdZZ66Ygpjd3/qwDujoIxkqveJ+d5jtugkbRJDkzH3rSMpB3ui
LNimpTzb+HWdXTCojcRNn9S+k/kdvVhUC50jPUMWcOJlhNHa/Rf1DN+u812hH9YQ+sXuY5inH8yn
KssuBgUA/fj4utGnVbad3FsG3yWs+TiBP7E2j82Ld7NuDhMYgk7lPEiA4g0coBsiHNYtWc/zlJRG
rVHGuT2MmRoMk2cBTqcTdY3LHlrOOGJT+EPiKZu7EDlv5/LKnp6zAZjJAehdQ9RPipwiufe0/zH5
dFHuXyGYEfKFSw9KihDoblkZQj82Qx9Hn3O76xHroEPgkiq7/9pU3u7LP/SeaEa6kGyQOvCtJYkt
q6Guhl7SeyvIbygGtlAf6uI0Sb06fwkpqmA0aaTr9DpkEG+BuSAMncjpPutw93ZubrZZqk0VOi1A
EOjEWPCE8z8wVy9U7PFjCGkkQqhufrjYA82W9WnF4ZVPu9twilDXlzRsbEzY1bnJPLcp8EZM4vvT
flpF2RU0VrHYHuvqnx+/tZgrBIEs5Vm65kqxmZ/Ihx2htlLvUSDhGHojFsai63G4j5M+nJNRshXs
tL4f1MD+kGhTKzWBOt2lPzqdnrl+tvnue9aS8JXEiMrUMZAQTfeYWXjzQKQ29FgLLyZNIABV9USH
DFbzplc1zc22TY6+rj4w5kiuHQVri6/gtRp1ObZZzJPhynkbmAE+soh5y2HdLkLy7aEYhvVsir3O
wJ1bs+pPW33qedbE+wC99X9UrnqOLUODBfrQjzG5Da1vW9j1P32OrHoaV1nRsPgwGugKHsxNjVQN
aik2Z21KjvNaYajIKvGR5ep3f5SE01RyLWwN6qtU+ZYbpTg0rPtrknt3Ax1niZZMru/WOnjntIU8
c3RwFYuYhTeuffYzmRC9dzPsI8F133f70P9IQceLytroNcLidG4C6JNb5N4oRSJm0FQ08un5R4nt
RUvBMBvNQNYnblvpUtngJRmIOXRuwzgqYkTp42KBaAH/PkbkZArWUYPO6FBhk0azVIbVW30uCxU6
neDrHYtF7Ix6aetiT3EIeFe7w0HQ9H7QDBQMOSpLpy2B6CjZuBcvbw1rGYFdrGoWnQDPdVF3PPT1
nZJzKcqyVRhejJVYXlrjK5NKeHUWdY2vwwUDwaIZ90jwlzjczrkwDXeUErKEFjDhgt1k8t6I14qd
LG5A4XlrXUh9dXfoiBaxWhCXFFDktjT3EIYF0C4SCkRa1evYqs3H3Jto5qDX8yOM9BRGvLrwf3Io
ljidr7xQAmMx8VKJAI4iUUjJ99XmePu33xXkCKtFQLxADLYomYM0shOjlAON7uQlaZeLGISXoHtM
FJ77ha5aOS00cKweX43qJJ9hE4TMbm+EDMr+IOdWRN5tIG5e9nRo76IyON1BkihrUY0l5GhSPSeh
wRyiNjrWOBVjoAcVLSZmPjVXmPsXQLHAo+HXqUdQb92GifiaqseSOI2X/sKc4Zzg+Xcry9LOS3Cr
GMWlZue8+spQjDgP96I3bz1Fm0MqIitPo98t5W1uTICQrILamZnGb47lK0E24UNYLkL+2ZGV4Qxm
Uz71SxB2wIJ8hZZh7EzYCvxhNLM5cQ9Xf16g5kn7O0uSGiEHKJHmHT12crBwciGAVkLuNiI/7k8U
39V5yDR5ka7qT5C/8jgSk1dcay1PQTdtY4SF3kb0SHq7JxAXV1SGhbOi1nNGt4IvFbJFIcsHMJdI
KyidLUNC/ymJJ97b82it/JAdJiuCDBFXAFf05n7BdIYfykkLU+jzABpyVhyv+NgxQixww7pheBVR
heGpspT7tc23pbEE5DGv6Xc9q37+mmY3S+pRDp0kPJAur4qMRlLSKsOooUzsWPuZng2XfI+ujKkv
2iervXYjjQ1I3sr9+dW8zeG6uZAnj1lTmDSpfTZYRjO2OXAJaP45LSn+0I9YjPAtGdavvtRBd690
g1zH03zAPYYJn2F738baoyJtFF1yIXsMWqacn7YvFAWkeLk7TeRiBQs3pbVSW3RfU0FlvS2XghKA
c6EMllNI8j0laigjkhwBoPNpViV3zM96dbTUHGRi9wTrt+rR/1vFpFRSpy4fUug8Ej+3RmESJwhf
oOCtrCFLPhWBdp5TlaeXvjnlb7dzeGwct4/yueL0UQqpfzx4g24TBoxIbYjGnqlrgSLfLl5nwtGL
IDwEttyyX8qjFwAnDqwJS/PSa4M9W1kaHnzyJ7i0KPzb8gQk9NV65awdmkzMw0q8gasNvJ5MFX3C
rxvcETSAqUXAccMR9MpJm21b2ZOf3Wr8TH2O/1Nn5xDTO6chAqCZyBf9XKYxEU3OxQPzplCle2Mq
Pl2ZJNxiQ57BRPVKCL1Jgm+StiosQF+yfqULBZchR5fUNL7vGVTLg/+V+u4DGhDuF140xs7XxETc
0Dr2e5D+VrpFlRiVHpKyM32kxQCGAch3hymtOmf3BvStrKfkyMs4brPfv8aoHnc24lFaD+0Qf2Gr
fd4GBu7ZisWBZiAKNgE1OHytKm+Yq6Oww/oFbaqieVYbCaFqa8bvDGpS3HlGjfU30J465TFj0UqG
2x34b1Te9AOpEpXHILo+ZyHHYQw8JmR5X4RvQRwTiVtJiI8NYLNo2RuD4SUAaLJ8CGTi87aZjBn4
tRzc9V/8LeyZD+0HAXKOrG+s8hYDYKl03jSODeGDXwYusxwSRiZy/yHa43jf3IG5LFwcOCF8oJp4
CvTN0dmu8yZaLEbpn9M074WGsaRpba7vlxGqATxu1pBOxo2Y/kjKVWA4GP1Kz/QQnQBiWOubWxoY
lFQcoxiTg7Wb+k66JMX/FWXxfhwYQS+baYQISbbJ+20/IZbNU86iYljWAZi3pFvZwD4tPKGQZb7C
rHEreZKCy7epi1m8aOeX7SjCjKSDf1q5l6v1BjeibSKkzY2abyfHr/i7QVidfDZOybCuaJru/ETk
BaATTCKORs5zepojQVi5rClDXkfQg3v9OZT2+9GZMt18nrcQUqQR1jkJ6bdQAtwb9IHF0vDC9Wjb
wD/l/GfGXzWs8OjiUVHFlcyig2Q/kODFxctmvPR0lNlGeVwPATQ50uL0LUbvaijEro5BnmPPiLt9
jBXhnzQZgnQXKHuC5fjcuw4706ZUG11xD/qX2QRPnH/dP4eSrZKETKtiCG0xqn8ETqsqfO+IIF+E
6LiRoZ4fN9KlYiPA3y1EQJZpCUb8eQ+ZbFZ616OATomH3uHn6T/I+qEZMhwLpUHIXO0q3pyrH6my
uJpnLzSyvJelaYgKF0w9zDJ+9jCWhM3PGB1+cJdl4ZuB1UeFgLUaNtgQPRlLgYjMi+tfn86xhvy4
E2yBft4QDIrlwvV7cGRJQfIp1fpIxGcIHhPcJuxPjTpU1JVubNNSzSNVY/txLRDRMpspOLOes02c
8/RJidLETOPIX9j867v6HR6zM3ZMRRRTVUZO2VRYqXsQIxVJMhURBKhec5G2qKAuTOUabE+RP1zy
XEYfJvi7wAfQCLnCLIZwZyFg7zIBQZ755WMK2ffy8G21HI6gjxopxkT4ynmrpK7W8RIkgL2/IiZY
gJIS4dlkGLIcXbHnvuotyTEERxe4x4mNllx0B9f5bpKFpV6F92ZR8jiglSu1QVUH110QBnqsyz0D
izb6qoEi2X+u359mz/rFQxb1VLVM7Hyha+zxqESeBHGtE+2VKpZl4LtKqNGo+7byqpp/eILAfZTr
FnQ+XSOAUcvHyUzPgit9ot24Bv1CPsZ8LkmtQ0jzVphOUjNm95m/kgLJWwve8suP2CsJcrlArvI4
NcYi76Ga85r6h81lz4mEDOUqLu2rcEUkA1Ukv/CH0T956uHIxrNUfHFcK/skJzM1Tn6LBDf5rt4q
CKaPXTtkalTDCenE0NwRWcUS46fiXBJaDmztjShGTA0jYFoGi26IyDMIN1WYdF3SQQ1HW4w/6BXm
0Q7Ewo7wKcnOcUWQMZORicI/5FLIuE1/cNmukHLTB67xbYSfBn/MzVK1bVBdhOUgLsIJQ37B0Fwu
xT9h5lSOvF7z5ik2eJXXsoCDJZP0c0/TY+dgFZZyGgEfSLlBfhWveczBkLMrHzIeHSYz+nYK1BRV
EuOYDRWr2rq56v3Mlbq5Ta4FsUznPJWIwnqGblkkwWpEyyCq3shLhlOYNdxygCMMJptlMe8StUZp
vQMD5n1bbmFiFclhC37HnYH1KdKmBzNdroVOyTnrHy+/Wea/6+SzKJceuHzR5OSk7l0ORJREgLTa
719frXeZklaiQ4b/Y57KTgLqVf+GCpYDSo2y4xq+6SfIccFbYkzUpu79oVM1nTAGYUudF3xSPh21
nhtOIY51msqrbY8abXL2SHqSLMCaHZnRD/SeTemN3e/UYQDwWX2l2no+FV3SCZgwqU3Yf0MHdubV
F5wVrCplLpAVCa5m7j6FEkTAaEbBo2occ76oF7mQy1db8LZvz1iDGRzFVoyFlAblL/HqfnaprJPo
eEaA499aIjUeYOV4zAE3lEAx9jjmeKmyYjr/Eh3Dk6zdNhWs9pMim608Oe96EnzvLA8mO5sODA2t
fMCbsl2D9MOj7Y3R2sYtkolWbvf/vj6CMvijvbSw5MHTn8qj21o4MviyDrU6TaMZKuBpK6lamXVd
1k5uiAwe8z4KaXKUV5+8j1jIOtqrodnZMrIQ32dSxMd3Myo5Tbz2Isz+BJy4v2tg9506o9XLFenS
Gi+wisfWmbENjcotBcGZ3P8l8yA5P0AhOUbuKysaFPbA6i3sR2DfIqLNiDajoTF3bfMtIthcaf7c
QrEq2UXpFdhboWwGR4qyDsLfBkmNLXWpvBi0OSeY1zT6hdJjy7RFbUOAKKWDjS6NRft6uzBSvbEH
GblzJpDbD+H0AHXJQbijY81zzWxS9IcqQj0k8Hke08XKG21ry7fUIww1s9WI4+9NyA6WXKel184o
HvBpswyRLJeRrKDErp1JmP2cbqJ8Suyf3gVvr5Z5RBMlpPOfULC3NZh3Jp4byxQmx8AcfZt+REKd
RXQPNauWPx+lYvIJAAoiqlFi/7OCQo+5d4aEDuakQ2BGRUJ0TOM3fdLWOZpsaf7L4UnWAxXucusN
Ry/U7IOym5tmJszMA2LUBQVK0qGrUiiFVPba4mD+sWZAZ/PRBjfx3sIiZbJLjg7RMKvhCwSL+rrX
/71nbIFTkxByUBqTfCb4VjQE2ql645JPzRTjRn+lg/9jneh6KahA4OdZ7R9Xf8eGTr6VLewzi+MP
QeH+HgRsWDAzN3RTyfVH0TDK+NShy7iOS9a1585C3wHvgALm2LbC5fP9G9rgflNu1K/pqpvP8jDl
c+LuwUxYLXX3iPNoN/2Cj2fx8Xy3fDnAoxOrpiomIuXE5CvawSYkeAPpVA/Pk1f0wnFzgP5DDwUV
VYd4/fC06ks/TcAHQkOUP09l0b3TMee4N5lXtwrjoQKt6eb66advH9vEXp0dBjTqmRlkc32Ef3zi
GP6d5M4N2NWF2EfTcpLwGcYNhOrgOnykH4A2SnzS542CqUSEwrTLmYm0cYuCaTRAPVClTS521ZRj
8TuHns+sunHYSJ4Nq7hhtkmZVqvwoismlwVl2R6e71IawMrNl84sLcl1vnyvOvym+4zRZPA0s5J+
lNsUKZE7lIOW+u4G5t//Uu0Earjd/jpRIda/3FgZr+sEfwAh5jqre0dLx3I/p22xfBvR/zr7oI0p
7g7muCOtqof9gaymqY1eSvCmFnVWl5N6DLIF+hPoR6VKw5Y+sHUCHs17eEE0UdVjnP5dA5peCoKK
Jr4zVVkvKzQEcLt1yHBELV6G2SzSsgmSLPklAk2lE+tghaaKqN5cPSmdZIFNlt35kLfaQUHEeAif
GbZkUJ2EbwxxI/jMvEi+gM+hjIXLp4l/sp5PRdikCzK1TgtpSzEuuvysX1AaWn5xn82GhoLpLXWi
OS3Dxg2tiTHDLGgjxgV1QedROvk1jRyi/klZ0PqPD6MV8T+1raZh2REi47f8b0GEqeBYZlNKgMnN
5hs0R7qqLc8v3U/oWU9afKcZ/zLuppvqSDW3P0qitrj7xio4mR98qmChyme7tvmjiwoHFBt3BQYs
pt9xRZFz03QosmoAQz8aNwSApyTnyphQok0hPWQjO1JhVIGhca/sd+k+HgSKD/XnYYNGRJVdrp0e
5WdUkFpint1FRVJ+JfuN1z90kdKevQ26t8DdEJFBavZgEu7yQ4VaBNOYCTqS0q/FnFOK77ykGDIf
R21j3DAfVskC3VtmSAHjivrHYUl7xWTpPaacb5WICDD9wkR7XVMGb2stgTwM33U263EU/CElr2Uo
YYO/bNB4S3sMZemKrkFXO0k1aEvSUo6SsLKUsnOCm5X0jw7/hG6q9vhzBk1ifESv96VIHvJxuJTR
YYLCUNYqe6KD6xiy73PYzOLZfAAqp0ZRbxtXTUhzqoK9EGVzhQoN6W0DcKkHyRu1JmGJFq5zf3/m
nwTQY2XmY785S/6ZKO1QbCfq38RpxvBgp22MRYKLErOZ1ik1VhrauFLIFTnUgTJ5TWiU3S3myAiV
eLftBxaOtZ+NbBraPc6xHgJCCb+R7YtDsLfAxFD3D/nCaKNAlNnthM1ik0cyZE3cv7tYJlCvpvd+
LhS4BBPgs6xY9p6mmFNDsXrGRETo8zXnXDDR1HuvoM7RNqqf0mNbzyno5swvER6aDE/YgJxUg1E4
ZzzshPPvRj/0miH/lGAr1RW4TooXIOjUhs8BrNh2Xu0890QzcFW5/uPzgAMAmLx9FM9429ezI1JB
wfLbzAPuq3cKVwVl4EM1ZKbZvTE3bPES8rTO35I6200goQW5++RZn5wowsUZbn3Z99kwx/cQHjMa
U0aYO6K46X+2CMYRV/rsN3XdTKLFgIdfsNqN4QU5tEmLEU8S7KDSqeQ36iYQ8noWt1Hb9P5f21jk
LEhkoxUtvCBNPXHIeV9pHcebe6a2ydxl0WKNWU86o78NkShs2WQ32W/0f4H323/4q4D+Tv8Zw2Ph
84yVg3x1Z6YfEMdoIidIFcE2kd6aZXV15zhSItT36GYl2JE1jFZQwSjITJYQJfL1iK7mutCVTJ8h
zpnOI8YxEmIPVV85FqNGGCGcgRCsIuglBXNAQRgP5X6YRTD7kL/pCdjb+1QPjYlzlaEJkJZOmYAQ
L6m59CUykmK7S7KSifSAxdJOabVmouuVE8qOLXSqoBD97eHIak8wK/dnLNbLmTjdu4Nh8UlwOr/w
btaS+pDl/Te1iWTaKjyjbAhFxClVy401lGR441FA299PJlc8JPbkEmGJ3BE6gl69glbK+mgmSDBJ
NgiaeZohkI0bFpnr1LrbbdMbT9aX8jAGK3xZNFMWNMPlejRXukG2LGz6IeEDdBW0180m4ruHPdQw
c5WpCSdUNQvONb6C4bwZMrYLyL1G0EoVPYkfY2XCUsRzPVlw0YHMkgso0bFc5ZtfOwjR5S7K1KVb
Ll92nIlo+5QvPakupVN2ypjviJy40VGix4yidOFNwm7/AVC41cOpAy+pGFji2TcHyOHQq028tZkw
Nis5HhEy6KsXOiRad4ByI76gsSIbPKxNRybcHnofkqmFyZkqlYmYGogmXxddgSDZcu7yMWAswcKn
OKfk0GV8oo1M/xuKQtxR/SUAbkUlf+JR7eEVIwgQcdSYmXUCIHQWGHFRqWTFkTcVW6JYi3XSRt6g
Ti2EPQJUT68DCJoh8rGvFtIoikNHzS5ZPMvWx3gV/FRob3cuoJLCiefvblK4/GgOj7TE/A/C2qpq
lyPUIoPcTCCYgOf0AdnXu95q/1aeh7c0fXG0RsnssHu43G/BWkCYq+GxTC9/7Vn8fROICyCg982j
Q29sTD06vol/pV8n0JWhD+Di+FTJ66wiYH0tksZPOkgiv9DOrHBWuHhFbnYukoCo8XBHbU9kuB/w
sIfk0OFU+mPkQhXDlqpWOqgy6/t+wIsnMAS3cnZN83246WFZ0csD0GVVBOFufi6FYeaaUZMYLye5
Nj8RSPm/sGFtBdQuswZQuKDlFS1hlZG4HmhNH+qwbkqtrCjzS/AUvCV0+NVMz36VOi+xEgtK58qy
eWCoi3VYimTEZpKVZjO0NW03zKenfabBCxsKmy80LZiC7zpUih+MUX7MP/Z9EZp4rlwY9Oj5maZp
iwu2si5bE8Eh37iB3u0yk5bHZZxQ6ZKhg1LJ6EbNae80irWTPeS1+l5qTrx6ninuEy+7YjitXt+D
/u9hCgCV8tm409NbjapFAKp0YFRRQBz6YjYhti1RNMOJFki8soExcJ3UxmNJ4ZUPmRkOPg0eVXi2
uLvliI7aicrI1ig+eFlFaheVHeI5mODxJwKbjuCTdOaYB1bygZf56XU4Gsaz34USpj5Q/5N9keeR
DQJRM8T3YHg11B9BvGdrg2VhRkupmSTwrZP2jFdg5HD1EuRs+rUEoEVaHolLjAyrgPpfEIxXGwsY
+vrISR08usrvPqSWtq45ISdSQdW8b2ow0d8T2E5dk1QXJV30ydHnyhvguUs1TfZW9owBZ1OGZfGi
2P/+dfqwhr+hHIv02t8NPo522DTNLca/BWXt1Vkbxk7IwNrPN610Q6HTxjvvSAuNNOEr8QtaeNE3
webIVnk3nTTcQCIG083Q4LQ4Sk8uJ63PW1qMqh9sNQvlgwaEKfUya0botZdGeWI6vbKVaOy5UcDH
uUOhvEpZrWZuCOw2o2HxoPcBMdUslbHnKSgrEDviZPWTnI1fU2uKKCtpdVUCYXpYj2td/HZ6CHBx
K3fMcolzEhd6IfPVyDqDJCoWmibmIP0wyBSwnDQH60mdS42VbsZZBsRC49qAeLrmoAlo2PPuu3b6
sFifiPhm0ZtkzFa01o3ArbYNsI0p/rEq7bOfEEM2znGPdWB07XcGJ3+9n6J513Jg969vMM5AHw8t
n7YHpL0g6817+XrwZCX7gcvgjtL5znN+cnVwH0ZBgnvtDr4PHZuxLfBCa/C/ZmtG52dFceEKvT2j
Ilw9FAHLtXtXu/XU93C0aak7/Vgf4/1hy21+o31xETSmjR3R5ydCwZHalauSQzrQaPbJpvgj4NRB
P7aGaxTRWpND8S9fiPJPfJAROSQI/vbVAHOqEfwQCuizCDokSaaGU9H4lKfRq7s6Nr+MnOOQpZ8k
oWnpJl5CjbPsBDKv4OGmlhyKTp1fB5EPS7DodmIq6LWihLmVYq4UECk+a1mfl42f4SL5wl+VZO5/
9TbKzT/YkUPY87PNr7XP8oIhoqYTk4LdO6/ribebUIbnW2bzq/CovR1pQYmx4KE7uyvZQkEkSe0Y
0VjH5pnhghM0lCtKCMmfYhSnbz3LGX1J5Mb8Q/blW8Rq7wzx8UwwXw9Ind7TnRjCvI1MUxwWSPF+
0EIlcNszfkIV+mkEfpsyZ6oLaEQsDY7bkE6z7zaBnzefetKdd0+I14jIO8CHxtKcBC4jqMwFtP+G
irPmWMX8sdPNYl0+CrbCNyBVe5i1Cu1V9pwL3fMQyHW6d1itgesRKxyFglk4atz82eBKtEw4K6Rn
1IewY0qWQKIi4mprethztd3hMRo5osqw1anc6mMkfVdqWBpJP1OYctTi4T6X3Z9FmaGqe2NkHCnY
tqtnTMPbQKj2fK/JgAQgASFTLtkU3SlYmyXQyimTG456mQGeQUzQAQl7OEsU+kLJDqpj2MV87XX+
+YLxjHUkgYZ8hAui8a1znRE9F61lFn+s0rhkCGj2A68ol8f1hU1P+6snYJDjOysLJmDRPqqPcsfm
MGqaJ5bCOhx5qfBM50RI9ztcHM0r+BcWnhGlV1SofWE2ymoTPn5ZsBy7Y+6miXu0QyLrh+L1mUUW
OnAK1CFVqpfcalECkZte71DoqRlmrqqmQagGaGDQrEbJScA8SUWdOX9D2tcdvcRFgzIs8w86YDfv
Q/50aNgrqwebrzMwktHSZyhmAFika1QGVjQTNx6+C187c2/RNZIcA8qpHGjf8YDVyWpZDA7qKNJ9
57e3VVrYAaH9OeoJAJ5Twqr5cYYvKvStmp4xr3kUqa+EzMVoG2WnXX4twhQOZUk3PHaLmuiqMO18
FpRmRHfEgLu6Ofb6f2HvL21gHS5EEZ3HlQjEFwRlgwTniGy1MmD5NtUG2/DAPgiv6orFlI+FeLZW
dzMfIUWE49RsmsOqCRKKQzV/pNE2JgOiZaaYuBIhMooKsRgy8m9TCkf9fZIlcHmAxoA5xEmjaQp9
P1hmNuQgxNpbRcTEV94opTcNwJBfbOjd3uKJInbTh8KiVuEwz0V8W25CcmfbCmS89GAa0xDD77lJ
IRB//FWEv4DAbhEUgn5ZLU6/hVo3oQ0BMEbPwkNwI5QUPFMhLSNHj2/ssKPHizJPwql7olRK97v6
rIBhF4Fb+46y6EZQ7x/TP0etSoODWno+3Uco8GIWLH4rYy0nmwy9X2RpMayYZZPibpj55cr+Z/E5
5Pxr6LUux6e3pEaMEGDnLMAIuN+6/XN80SZTuvlrvfMI0RjpxrVIxX6BmjRtCl6/WafmgpzeiOgY
TNSWMMlgBLSQ1XG/2SiIVpbfZzoGphHDA228zLK3YXTYSs1LLsKxmtIe+Zg4//hZNkaRB8bqx3Z3
rOqOtiZMqRjclIThJhcYUsfqQ0s301g9/WOYJSViIXVGoPvg6iwZROnSZTgvupC6m1c848MxgPCq
csMjskz7jgiXwB2I2Lixqm5kQOgNyrZUGywhn/BvXQ8d19V0jQxQA+8tDgoMMm9QdRoRnmU0IRdf
s2h5Dd5pxFzbkwxzGH1XxBRzjYwPfKD5zPWgDPSZ8Tehdl8CvSeb4M3bO28p/HKUjORbzayhpNUu
rYxs+0twqP7/shFBDshLmltvu91Zb7u145RMgbUR6GGVpwrIqD20e0Ow79WPu6LCNrI7+5/W79cM
74KavHSjGt44ZsmOyQdMWM3OuNIYX7S4fPQxl+LVGRfAcHdxGfAzFaCAODN6F9tcrdATdQBnG5yb
z8LdlVr45AOdWu1QIqRkMaY+uGZLUn3HiNYT3mbuUpqbVl/k1YCdD5tPXgdBvWKCiRO3BJcPQ0iz
XKYN7moJkzgf7DYYCHDe8eyZjPYSXk4LmbdOITxQ675SrJy1rDCUTsjw+MBnseaWiESxX20gbRbe
60oodHJ/dwPMNr9uagSe9BEG+/kzFY1rd2M0pHRzFX2NeWmXHX/lqN5UpMoj7OovF2kREvb19EDd
gNunvoKHE1UzEPxG4BcB+uYaJFhRQqtRG0Z4//dGloES7+KSBm5A4AU1AxhGSEErt0JuoWWKoeT0
9Cog4PFeuYsUIlKdgEcyB8sdlPpSdJO1jXDuzuFhmRehQexaS559V0YNCU2kV0/nhF022Lczx7h0
DdB36NhZD/44HieJPrG1e0HCAxX6zKoYVD3oENt9vY4WFizlnCel6qxeqPlsA2jFAH82gXoFx6QR
+wNJhPWzRulaXjuG7NptFXAqn9MPWhlBIuExFTWbSezLBpFWAeah65YAqxGT55c0/pWcTjI50dqW
fBY0hW2mGzWIfCJNdBo/iCM56sf4wRVtBvc63YcYOwSdrRfEJ36t1+7sAeUYuaNOhGWmkExqFWIq
93aYjZcC7/qql/SKwZcbbQMOrjGBX2+02ZtEaWI5a9L3xX2o8CbbTtN2HevKX6CoOkXe1H3Jye4D
Ui+lz6K1QkQmkM8jSYXLACM6JERI8OeRvrYaiLT3BZmoD321PkgLUUGi66DtenM+xVd3rLf6oTgF
4frnvSlTMpnOqds4kVFD2hznlDNhYYspZ+ngFNmFbWS1cNQA6bsL3xycLBw9xUUU7/gVO9WXkhpP
KfZO6qLDT5poGwKioSEVggma3EbLoerr7bX6BbqGMm7sHSlaUzWbFHSpw8TFNE03J9SKfqTVNDYu
3wpWeX6mIRYIQbTncEHRHUNb6T4tVMUhaKS4lF5WYhNPu3JDCAimfkFk11bvGADm0mGvjIWTXh+T
sUfXyYkdbyD678ubt68vkvg85ALKyzjBAzjeFF8AMHoueHLRnbNBZ9UfKHpP6vmUHIDvqMByFW18
OXGaaap0gpjqXuyXwdigF1WyuoWNc22gQtD+yoZTLClJFzbQ02kfW5SiiV76/+nRa92SOS8QvXIi
LAanLBNmVIS7Fz4ZSgLPa2EWdrrflecDfaIGv75UHtBMCJK91jdsbgGdD7+cwbSkymWeZ1Fu0056
hDO4IuNJQv89335Fatlgzq5GTy16zXPBkCWoCbxM+9VICs1OpaDl1yGve9pYIByFYW3TBqzNQacx
nY/zDHZDb142OXreqfL5R9cUtQVGeIemWiSboJRGvY/0K7q0fVb8Ramo+8ZA8j5UOjW8ofsJIUel
y6FW7aqZNS8SHbZc7rRazk8HH1if9eaqZRKHg+PukX6vjZqglPUX+bPgZ9Uz9tORS9iYRMo/lxXg
A2iPWGJcbL2RIy2Kb6l2MRRwbz9TFDn3xqz7fT5geAfD8UtFRTKHRspNKWyJsv8CGeuHPS6J2nbW
VS4vkHLmdHWGSAyubrhhGVVsIT3x618Qhfn34Kqj3W3XWRcfZxZ+aq3PNi396HezWBJ51K54Qg+D
dcVZq9vqOKOhThwEEe3BCd2drOnhJtomIxPgcG5RTVIB2nEn2LXnXhgKUDQM/cB/5AWu6WYWepGP
naq5kJOS7rIwtIhaoPNFr+TDJ7+j0PEuUcGuSR7n5VMQ6s4oyLfYQujC4RErNCE5gh9B7yTxFWkT
TCWhTPxrrpaD4rbP9juqEnbcC4UQHjVU1A+cWJVCI1u7Wvt0ZObkcArMFt7HVNVuE76Z6j3r2LXd
PhM9GNVCmo/tp2l6WWFPlNn3qQi5cEnEoJTVXIhuKxilqjEYtdblbLU6qsHGO72K24RT7VrRkgne
sF+6pD2aTXvpQEvwMxSuuFQcZN2fOIPKcNFAYKindgUlqaz5RtmqloRd7aBq/uZ0guPhc1JuIRLc
HYiRwONAS/HPKH0SDTimy2bjBjX/jTBWlqSypc8Ppg+NozdJF64GYdAzROJd44Wb/xBK7PwQbIlM
V5M0gjVY2Eh+jr9bsjDBTz5Gv+dUWu6rbrG+eaEhmDRWYS9E0BWWiN0+urthbChWeU1j0dqHBsuY
RutFwR5kaj1XS8jrElhD7acZpVhq0kxVbKLQzBEDoAMSQ9MOgVKzB+w/dTNjgxBHqoAiYCk1bpyn
GdsRMJpJwURbXhX4s3o2KT3AlUgnWD1C0e8UtkEIF8q/qtnu5prtH1G2lu4dmbHRlstyvNFbtwAD
NNtPiu9yk6WRwHb4CZPNOejpoAiOFRihA+6KAhjZB6qhfyMbQJUwi1lS5uZG9pbQIyKKT+FWf3YH
ANLjiGbx+9vp8RHQBXb2pdDEZTEJAr/SaToArGIGZhloFRZYXFB9GNhk14u52j6bim/tibJVUttO
C52xgzNXObOOiDVXTrqRiofebZhFM68uMD8DIRFFbNhOE1XXzz3cLxIwED0pFPUBS8cAK2dbH1pI
Pe/lgoh2Bz5H6oJQGkGUF+QymSL1A9W1PlUyhz5TleSbFSO80u+QFaiAnoKr96RQ6A5HRvP3Esfl
COJznKp5wuxo804fUhoOZxXjAYRpSc+/yhdp3eVr3aeNhw7m4dmRaWvgbMrhH2oON3Bfr21k4eoa
YfjvTM41sEOjX8xdWbXAAiotf+3TWnlMrhIGVgEJ5RHKzf+tKphBJbazSiTw98HszE1qOt+Sd0T7
zxaimAG435PXVm0QVxYwgfs+NpGPPrY6tw/MM5yJGBZmH58Q197L+DpL+tTd2BnPnvzxYpDbgak7
a1n8mVU4jnD7gC6ZGdqV+1v7fCaQsRfwM0woOSQIzPZ+XOUfKbFPObR53roRP0ruqxktyM5dJp7u
SVDN2VXFPnbkkcQgk/+cp2ufj51zPEPuFBmOj3T3kUYG7Mwrq3OTNgsvmINAnLW2WntaisWBR3hX
mG7viWc5dHGyl+fbH1voa9bs5Mc7PWAqYCLgkRzVWfACpx5U1PSo4aXf8lqEt8DpDfDpy5A4SvOl
ZftI2/6fwOejqinpvD7HYhuZAImJD9cgyC9vbhItXHZyFv94bstB9n3fSsoIfCLcXF/TO8+l1lTC
i29Bd8vtybwLS80SgXEIHkKGGNJ7sgPSS1B2U/EKb3KogeRwD4GQFgG1xO++k4J7i6kah25oUW/y
T2ig/VOsaYtvHp/DXH0G17AZQhTq8//rha/fFIxbu22pQd6QxhRLbCM+0c5oQnbbZeR8uQ90ySma
D8L6I9kY/KSUxGqDbvj6IqSB61gPDN2n+fmM+Yzglb4dpCsEUOsWc86eWnxJiZarT6R6s5hy3UoK
687/+0b/8XtxY7vKcNTkLFBeNzGZ2KpDFqijBr8+NxG7lFmd0ltjvqnZbebgdBUHkqwm/r3NhmSN
VE3/urFzsYa4Gw3K+qqIEkJItEhYNlh2ZQ5utVHF7yj2GlOJGs2SF1DNWI6fU+uSO6d5m3Qf8r1U
06L++h5EYn3/XVF7GuxKvDxFf+OQYy4W8xrcPPaSV4RCFLtdfihVhhJEQ19EZj6TtiZhc34Ad30d
vMr/PYInqFUyEt/ad/bis2z9gZz+cS6UV9UoYbK9rLiwbIV9jDZg0F5kAntaJBEoPqwlvSL2mZAt
N53w71uctuBklEC/h+Z9+sH1jETJaPeMAKW7S7PnRWnpFGp8SdCAFqN1DzHJJZ2lQAdSdJiidI7W
blxis0FdUtzXVTeR2cWhXpZ2774lIpDGROWfYYFH8Iahic/nvBm/8wdBhk0cfqm1Yb+XBRDlntqV
50pjhKPKmubvx9VtQAVVdGaBDKzHkjsBmi5fNPBL80Jbopy/H9Ah2zWfm/+XRHPUs+G32BNlnuv5
D+wzQbstQv139DilvXqTutsx3DkD2vMVjz9p8dmus5h4Cx4Jbq/wX+dkzk2YdM/CITEVsnTZceJP
tEH3yA0GGMabwOGVuYjvP6UMQr1P82nYOyA0lCIpZ5N86hIeHKf+qkQiDGSYweZIr1MTiSne2jy9
Es1xhj4Y6gBd5eZkdLjVWCgFKzyRXqGSA4lBSSKdgQromdRwjrJMjj8NmL5qk3DRQ91eMyZvUNMA
Sv2ieCruDR4/yCjkPNhMXY+C2EM11nepOSiBL9ItKsF70O46OAY39R0W+mA3l2V0cjnvqRhcfKoS
nJ3HiPytvdjyemXfY1Q3+q7lF1Pe308WeRf7xuB/UXRsoYkLlGw8oopj3PtyNlPjti2tBDcyt6N+
JY59+3Mv8fET6FFh9KYS1U3d/bTBcnhKbs6EaqxZQvzOMD31dyxCzA308zz85Da3+/f1hZIUNKGp
TG3HRwR3ZXR8qxf9VpXr0Zgd1+mDAoi1C8MpRpoKuoFd2XCn0eZ+wuLGKhSCyUAbliEwNV55J5VN
8TSfVCNq1f5kcHEJeBpCXmmigOr5FQBHtiWMJInGHlk73/iTFo8FbzRL1nXAgZtgfaPHWsbdAhlc
1sLkKY54W0xooVAZsdDNnOp+5ds3PVm/fdY+I8U7h7BOqkxEAt9Tr6Oy4mTmQ4sM1ONhp+DRfxim
PdDJXkhKcsQqOWpmoentE5hpyBWdrdqIZB0om+SxmUdwzQfkxsz4lz3MGyvSem3nz8f+pzGNwp+L
7fZLeYqf+mss7mx93qzbQwz/xoitnXbLSrashNX1ZCl9j/zDQt+F14QUHNjq7P6R9zEm/QB2aguH
l7VOEx20s5zYUkKYeBagfb1A4lJF7Roe1V4rPPQR0vhorLyrTx5HHHuqKp9joXPGVtQjfKomhDg7
sgmhBlUFc08Z1jPTQcgCvdialwUQAoKtXj8bkgf2IAUaNGqcpKe8x1MJomUmrBSklA2wTqlPNYjy
ZzECsxrhX1R70ml+9MmajN93bJDbl7TeqJB+Q3xWc5+hMc8e2xeNXzilWU4JdcDE/ys1p1W9a2BY
phmcq2yfU1qXLdo8bo2N8K33ExCHHhsP1OUHpvGr9UJs+hP75mRMwjZL6Tjk1qNZ6z3QhledXhqU
iJsbGpxeunzyMEnXOOu5U9cLSwMPOz3DRP2a3erbXrjuk8FR2eb0xpUwVK5PrBgqYk20eMy9suOt
MW8FUUEK541WyCw6Cje46OPApbEWQV9nAdaGBoa4Bq6UJRyY4mOdPILZIIU5SuRpEBr8HGC7WYa6
4I5+AZGJ1aUC8yv1/TVALoqFhCBv2xw+iiqVUrJtUKXlmhZYusETxo3fIIA+CLMw/bVBhBBERho9
TWZ8RTbx3tfpHeqm56Ptc7zS8dWTMxVCAylHlfwQu0A25Fxt76T7TgM+Dm94r8+wjuan51461f5R
PWP1IByMP1QfzSu3tm04zyVuJOnQGZsPW5rDOyxP7f6Fh3HIaOEhtI9rJAdDu3JbmLPl/t0uMv81
K56Bkh9z5gkk6OgI3kOcUedTUBzHRDZ9nwI41JqwMZW1aaYwYdfkU8YQbV6m3h90YK5j5KaS5zYr
WxqTRU3Dz/KqTjMQaHlWr7b8nZUMnEpE7RWeD8lCZsPbNFD9QtSMmOcL08Usb8QM8kpDFhlezvQN
+MBSE4P6CnILFF7u2+V5D18cDw1IlqT9ES3WzIqQ0tjyiEkBscAA8PBVThYqnOV/SRNQP8Aq0iGH
ZyljH1hYo02t+gUNU2xbKCEnfw5x/aielf2WhnawcUPibTs42iMCx5DgzFTycGs09oaO6TecvH26
xFfoCC1W6FHEEAX3aPfEfR6gmQq+B1H/DOdlDO8m6RMnFrNeux4cPz91EZ3lqkBPsYbmFUP04IZV
PulhyBlg/Rg/11aVMF5cK5mi8PJGZaI9idn0zktOerTZzlpF5AEShfHv3mRy223tTzAf4+ARhXAS
t8NDkFnN9bc9FUii6rBWZIdP3C6VqOVfIM5D88g46zu/fU7O06jvmf9Kl2A/lyLAA0MSDDjaRHBu
Oa9+a/qqKtebJxMWDow2uuY8hRlSu4uMO/Dorx/lY1WUo7pWpozSGa+lfuYReNu6eJiRZ4SKdUt+
8wIVhzmH/WrO45eolGgbDvhgzGSPt81PKHOvH3QnYhgDYgEXqNisH92K1jXQYPcrAE8qXNXc/1ed
gLiAtRoq3ddr/g8hiFj0BOiBcXnwSnLvfscskXSg/f5KhnZIhlnwlsMnXtGeHqmlC3MLPP2EWDaR
HntwwlbsUHsO4mKG/Bd4qQg0eO1lqOvB06RJJaK488GzPxPB1q13BtcZ8/L8E6HgpkVobvKfRS1P
hJGUQf17rQOnhZYkUTNVuDodlHHW/jZ8up+tFzSI0yWL7ccXgCmFgGM9VpETP6zQIz6tomc+pJ2i
cP5rlVs2DgAJ2sFUtWt6sf8wSHBLzK8bq/6mkTSSFPSF8SZaMrMfNECLZa3dbJH8Q/BHV05AeCQd
ls5ZMh2ytpCwEbFDCbfDLG94qmgJcGxrGgjDY+8taNiB2K0A/GFcfWmJ+6lMfCDOk2RxDaFqDcDi
dIGZe3EkYGheS9i4+erjC5AU/k4SqBqe2aHmsMZK8HW1APMZKlC25PW0cgVnmKOi9xUD6xVRSH+c
InAp9Dbx1y1X/Pyw/Lq8VSVXEs4rsWGJzaE7HbMH1mmE7mPbJB939QIgBavYR2cEuP+TMYNxGGe1
0v2hwulRTQMeTXupo1HRETJ1YFNdy+can3rcqVm65FiKsd7eKs3gnvSVuwkwjq0k/RKfUhhRJuj0
u6hNDNxYMe7Q0nKQBg6qJUxnrflwJDKmZ/bkDBCyjHX8zZT15eJ5lnt2WMCW+oU0leyuMV/7cJ2J
+3g2nbXp7NxHbuXnGQhbIoSBCPOy/7aT3ZhNU1rM/5IzvLkcArqtvHdECfwBFVbD0vt42jVaBu0+
lUH4iNuyl5qOlVJ9Dh316M6CWHW3PTyYg+qu+5zUnKAZIEr+rTuAlZUtguuCAHIP0JZIBVkTVJYm
eezPIr4UKjR980EO1m58MLtr7M9x+1CgAHfXWs1HGZXUACMmHtHCDf/4+pwBuI4H//PUn7EghHQH
FH9JS4gmtakW+5ZEARl6AxA9jXvo0k6nessxQdKGKfZDZF95VnCk3UPMHYZZJ2UP2JJ3Qnny/v23
WJsYoANODyY9iZZ97yhjSPlbg5K7YYXlyqtW9aqbWjWcHCzwB4Rl1TXGc+SEq4rXHiabbVJt/Bb5
6vOGZcJmCv7QM7fBf2t1UaR9L13d8z2H2Mx022OkjbqjJeRq24HaBE5jL6P40HK9mb5r/lDZhocT
f8gXmfEhfXO6SCoFsywaSSL1M8VcCF/T/UF1p2niJ96xPAdrwU3h39hvl7dT0riqVJNvXhYQ3/hN
BylDG+5Ps7NPvRMd9nSpLxvK/fep+CZKjhuD0b0kpvY09qShMrUIof7aRryonudZCXr+QYNuvj73
pb0fzcG8rCVrmV/Q90JwFgOmlvHc1CIlcrW/MvdRrU3DuwVLavf8z5GqlaNDSgAnkmo/rr6jEXGR
WpTuUxV6nKnV5LN7a1PPdv2z5gMtbFkkJGOxXoVVab4u5ukYdEhV6dQa2UAE+v8hP/gSB1hY8qt4
ADgmlSundODq+MrgUGD6eUS+0fvozbVfX5yj5rbZummRvC/rCdwfm8lgIIQCxlUeUsh9R5T7Qt33
LYq92Liz1UYE9nhWnjgnFmuICtAFROaWgZVSfJey3uh8pnx1KSxaBOs837jdUp9C30FmcHyd0uZ/
BeyFtDR1BafCSAI23ulpw8ErMiP30sBlGXMvZk0lb+qi32t/8KBuTRuh6QQ/mK9JEedtvQsjBm8m
qeyg6kYfVid3L3RBQJ7zhFCKINYKm014fwf0+bSragmftFgCFPVpEGZmXnKE8YHlUFOxCvwJwagZ
qHtLzOgJq8VOXo6zhpZG3uIzXY0yNr6+mQVNdn9F0iVgB5yISiIGpw+kfeSVZGiPuS35S5ERyzgd
+qMIn7U50YOrcSAbacEfHFGYNX57lVg/yjUyEfB+fKE7kspE0xwREY8xmENoAMvzDzVVVHSZLNgB
s4aVHjC4C8n8uYOFKj9B5qnsbkUN1wSSBE8WaHYg/z2mkwE8ZNaAa643+WWbUq1dQ7UxdD+IBCjQ
o+P8DGYSSa5H5M33uBX+3oadPCuZSVNR6KBQWhvzYj12mxz5rG52mHq2sYQn1tfXTAZpqGZRs3dF
yN2AgFwbEBOxLsEwg0M8HPiv+Tul4mMaePmneORyO+PNCQ4p49NasGyUkzVXQuvPOO+XjT+XSOtD
udIXNLxbnqLmNfT/nxRpab5FxBNSgzy3XuVkyfPIjWhur23pm/IiC2yPXloz+ifu74kJIOeoVzgp
TeFtttLlVDuHlD3guBmi3loZjDC1bO9fNsCn6U17ktiCCy2ATsUIkDdXBp0PWk7q/gMDLCsCtlt1
BOwYUJguOGIRTcuaf1UpMP97YeIPajUWcOUEwj4r4s3CU3+x491vwxMBcqEsN1RJhTg7fMYTKM6z
31FyDPvEIpSuCxiaNF38oGfW6unZfC8SxzzDkUY7xIzDrqCO0Z6KCQmzAnXso0SqJI+kJkht9HEb
NYT9K3cWS+i/XTuK2qg590njoObengA9uucynNXHYItA0Ey1gcNtKmcpSVZZ8KhjsUr3UnXhSEcn
qUEojzpUNhHj+tfgP2Vj+2L7uWXzFUAZsL1z3vPKk4N++EZ74VSFzZQwPjpT7gadgHQuz1mz8PPW
szzK7Fyq7CTvmSEE1dqN+VxeRL4GcDH4JpQi96CGElghNarJhGFCbNSyYbg7o4c3hrpMnextHJoI
cKXri2gr0mIOyaLrYLvabdm5qm+Ou25c35aSMF72E6Nh8bwE0ZOAd5V7W3y4fUOb5Wipjbv3tsY8
CKagiqMVKqo9GdHJfbs2QMu6y3zZGPMLY+MAADFwMsDaTXSeeDUERdnovojSsRi8NzRNzbEpbl4H
CgTMB+hlZTpiRG8gAifmTc/s48XDALrn5U8Jgo3FlMG9WWL6klmwmbKmJytYUMn5UEQKspGAWqF1
4TSyGYzj7QmdIG4klN2hT/2Gc7oxFSBbt5iVSxpAkM8YlM6IGjIGDww3euX3jrIP7lPPIVDXznC+
4QCro26D+3rOprSVJB6roFTe0eVO5UD3J9At0OAIaMzFXmqBJpI86ESY4fGwMablYxxG2b+mco1x
JNUz72EiWWxX8wrgVEIzZ+aHiqHKx9/P3C0xzXkXGly7ly+yKsvdeHoriCp5OdTKmjHJgk44/DbE
LGewqIiOXVVFWLsWSuahD87LUeiypMYU+ZduKOON4SuT3ewYfwf0oSgt0tjYGc3CFHVhveLSlIyH
558yxAjrXlV/1ipwBn8u6gOsK9tmIDT9uaWkbhTjVNVMKY0geayV660+t77hUcaY4hWh/NjiOA/v
lVEqV+SCbG3b6t/11uNLCDf06WR1JjqW9AEe9WRNXsnj/Cz4RNSXiVL2Iy6caTIP2Q/vEOwUBKoN
+u0qTBfjC2rqEcXdP+ZYIAcJKLFoNhvUtQKFhhdntP7UlRqg5FeSmOkW/E1cso1+PXwfuEATFFo7
sNUvNRgTTpzzhx8b5S/hmTnb/3ix+pSVPzVUzhqNevO8Vmb9fGK6YeMgGXiZDdzztZhUj/+lIzOb
qgRrMpAijlTe0KElYJ0Zj6muqd2mjiNc+Y+ILIJuSG7cOuoplfHo0gCfLZsCPQjTcjczzkDhJZ8+
RM7fxDveFbLg/0amsBOFRMCG27OVlevLzwX8pxLg9almfvm8spw3kdw1K9lYPOUZu6nicsXshsQj
lSSerMa0qrC2zXM2VG2yUu9cJgIOHVUp3sjoORNbDYEHFmspNjPZU8GAc/rqtVDVE2Vo0hPSWjKU
scGrz5SJDmSHpwT7jk3xbIehKQVR4bnDDM2NgeRvdG8+0KqXz7yatIoIGFGwBghdxxNK3SgxShcz
LbuyzwfVV55wYzIMOp2/WMxoxUrKLTghJntIixoHxeE2vAZcrBsZDQOiK0cifZqGsmHuHdW+WgY+
u7GgzpxJ1H7if/ly/O2YKV7dAdvdqy2wviLTk9Xboqg1U2paX71oY0FkmOGAecy82UTny7cbpuof
CLNvcGMOZh2ZvP4YZnPOKBNJrTRknGotqFqCje8C4hT0NMWorpTidGzUzv5Fnqye3S09No+lPoMM
ux4hrt9N4xujiSXT9WbSzHKtLDA3CWMk5mEWSer8RZaU06wQJIji3GumOIcT0K+jvmsdD4JPQC9J
x0WINhqoyAxDmo3UPdFvDONfB+d3Ut1TxouIts3AMRn8F1bibXeQ3HshZA/Dqk1ZVu/1AyED4OLb
tg82DizC1lsCPgRxGu+LFSPGDCLEsDaEgR5emIYXwaQwqJmo7MVW6cciRnnpZ5b5IUUTFDtSXULa
5pAMANdYSVLBFeRJKSRwNFIb8M49eBsOYqIbVuIDs6zFrXgriECIongaHsiMmvki2lPTb6UIgJV6
mdWb6bZqbEsikh7b4/BbxPFFL5+4p8xOgkPviSHbuGEDc+jbWfa+2+mcQanVHFBX9HfbSYpST1aT
dxOqaUMl7DATzbaG6Fmd8VplcgRFPI04mo0CZKW4QbYGop7QV2iuB2Y/tA4mWIrJ0q79gWzB2e+O
GwVOi2GMz5k8ELm0tpz8DqsUicgnWcJSL0OepcW8E79m+L6GhuFVcyw4wvYGsjwJOT812+2G/ncP
7MrvN+0xjAHibUUMf+CBBIxrmvsdEAWXmuDZ1l4HE6bdAMmgRf4iSGas0viGddv+DHcSzoQKyuW2
1llQDiM5DDD/tdshLipfHYrWbwKEpJOX+2msF9KEWfqxheoWg+ZIwEVOuKQPSnDNrU8kS4gMIQpn
fqikra6n8uoJhTVjeAqz6PDnZZGUddVttNoVzlE7YxRA/YgJ8s//1c8r6sBkXUgpAtuT7PSIYnBS
T1XlSE9o1APYA0Yz4Gc7xl81QfGj1XlXpG68YHj3Z+QvDRDoEAIjvNjKNDCMwz+GjZ+SdlM10AtS
37RZdk03HKbNpsOzguRjIHw2Ax9IlNIjZtmf51N/vhlRRV9M8Myq+kDlupnVbHNTsfMeVYM+z/ij
4QN3+gc+nHAHuqMoP/pLPjcZmg3aEaPLDEuAjZBLdNXZRfwpu6W3q+Mx2qxl8+SnRThvsEcYNmMu
Uae2qGOZ9zlvxWu6i7TxyI1s3e8mvl5V2IIXUrNsxuO7KP69AJIDHZm1cQim4/RoKhWZvLuNxZUi
SilcpSyPU9kwXBcxRY7UaGWkEOyC32Su5ZNC51GFvuh83I8KlcPpJl68QQkJHhFfIN3AST4mOwKf
tCBtsOVJH8ByfWBYLV+1PoPT9GpgNT8OrD/92yB+GUSvINh5wNCIF2AjT/YKGgDuiuSYxC//3Gr2
tQyBZODkfrzSR4hciRxkjGTE/4FwpuRqpapFrYkH/oEPwB7e21AMkRyXZOSg6l4uLOVnDAWvnT4u
74fe5wagtsJZZukU3ziT4QWoV/qlZXI9thBjb4qY277ahucJhTZy+tQi69o7AEntwBNh3A0fFEl1
Ply/aFaS7rlBi97a5VM3qY3taVrd9DlkPs629w0vzdK9KrfHtR+iHNdkyyk4CsKdUngP2oPzLaW5
H+A/1T8IgwXagq8XisupnF3Kq3uKHMiRuUTA2oceEU6a5nITiNCuimtN7Tl8YvEjEaF16ixS2lVd
fzMbBXSCB+FyLPS5xxSN8VfE3z1uxvwBRuXy3eJX+RONrdq6UB+nN5vJjOcV4vD9m0QIoBaAw0pP
H1Lp2RXQEiwpYCkIJRPl/WBywi9UB6xukdyDU+wIpgTBvOud+ecowYTcXq8slePykrlciFIBdhhk
BrLRCqJvLOItTXM4YUdUgI/myx41njexs28Smp0Ij3lPG1RF//rYugLgb0IkwFoBIes/nzFqVTKF
gWwKdhCYaZNnwl/Qp4GF3HmrJWapyRR/2LIZxNivXEF3ZtZvAShbool2ZcVj32LtABMxVwePu5Y8
YX3HEae7Q/aWnuj6r1D8nmIjENOxDTXdqiXrB61F0S80SESUoagNoMDPmagcSz5MWk86iOOfBHVL
DfaJJL6OVtsOj1PiaXSK8qXXh9G8LQsX28kXNJ4SZ1Mlk2o5EH6wNTnCmw27IM0HHl519QUCg7wq
6dGHsUAJjpuzgzezx9aVK6OyyiiGt0s/BXgaxZGsO1Mfl9825P6yH46SBDK+WJmjFNgXbvxvCd4O
IYtsrPb+V8wdzX0P8UsfiaLpqWcGcDCZTja0KPu+vmGcrPvW5cKOZwDlJfLljPZVMhgtebVt4+TX
pZRXFW6mDlanNZM0pmsP73Yjchpsp52zfizpnaJS3ZMU5ODLAZWMdcV8+I9/znYnMz0mzbGlE06g
xMo10v7DBwIHxARAD7gcuBmFoSEJP+TKyrqa88ag0UIAG1GYB7dKr8j9bJLwnxywMfMa1GfYywO4
liV7oet8v8+ufrsYz08jtoae5/AqvM9CDgLyPDS27I6+f2b2FtFHPGeJsDZ7XmNTdeWa6Os43CbW
Z32BkqHuSNcQyQVFbrLM12Eb5g2CdkJ1lg+sky45VV65gDrJUW3KpNkxDBAPCEbJMpO6VfoIkJwJ
jJpTXzTD7b2STLE99b46XuYjc+iOoaZoY3nczheCzyeGe2gD20O8X/N5dehTQ48emBqH7Zw6vCoL
3wEgr6LZW5LBFOybjTKgYK0jYNRjdI5FoqfVxGbwUit13mUH8Z2jVsc7R29oJ1chHHo/VX8i5faj
rhHnW//YY+rzcTEhYy1+YsajJhEjxf3liCoiwTHRM2Omb5eKmtGF+5YIvEEXbjbV7l6KZl3yD2aA
oofJco5r750SnC3KzFxpDAO9EvOy1W2HNSEAU+lhBNmd4BJx+X+D9M/MKhgizFM5IQUSzq0OkV+d
rQ22ZtoFhWqnZW2CUwM1maGwu7OHc+FvUOCpZsTRtDKp4bprpLZqcAWriOdQPjrDN1z0OqhBxe/V
xN4KZPAESzg43RmDORpkGShErilJ+o4KQI+b9o0YC1k0bMwJahwDT/j1+PcS9AJ2B36Lp/KRNWhF
OZ4S1YW54+g6HPZ5sbpcphwkbMdX1YC1qzrs3/Ps0RET/8x/KgqQc9/q3ZGTLdsFp0oIQEPwTiBM
Zg+bmaCVmgqL0bgZ7MjGtqoyFzAFm7ERaBejayuRGaf/fUJJHPjlobISPc9X4AiFyDN8pJ9WT4O7
MoKD5omTdHJvXNGfKb6cYJQUUYbCCVJA5lurbsuzgB+nkiHTv+SaRbNrgTfWxIfl44tL6pbID0bK
k0VzXIeqRsWsio/O8NpA1i3Ufw2PXppVPruDdwaPDN3yF/8N7YEjzL8uWQwWK9omzycdKNa1+QbG
LzEE05wSuM9LKgt5tCNnJLehS+oHyTFYuJL9YiBcJvdN87xrbySdcwMpv4hFDhS1cpuFbm7hrVA9
9Q8kRP4ubQSlyGheWAFmadbhq9Ue5jBpvT+PSamCvwDkSs865IHFMplzJz66NG1/st4jWl387HUx
efDJ91bdsacTuAqU0FbDjkIVwREAgvavSnWSO3hz+zj0dulN6A9drFNTEmNHWfvxg/EV5VPmicef
zNjg0EcMcLGynQxTNpyTM3KeAt0yc57Vyo5GXyKL7OozlfvTRJJT96qt4By9ns7gBO0rbxO/MJ0y
uZMi1N1Nf/0KLXXGaCZQdiVd85Fap46MTtHrXeZgjYIvwHVGBDGo/QMx2l/h7Q4Lllv0IymzTr7F
NXbIfeKwAXGlBSZIsMA83nxp5NvjOWXq8VuGUTaMypEP+vq22qMUAOnVsDNpQUj7CIN+TA/sRcNJ
3vAiWsIWkGmGwTfxZh76ARE/oT6dIqbDoqNLnCLvSwBKsTzGZBPtNa9yppLb6G3Qb5fgWkM0X0OK
btaYsggWm4Djm4lgkYTNc6Yw6NupaetPBpKsfu/7rDCVSNoZ2ii49a760rOlCXwvLjdUgM3UdrR2
HpENugzQwnmTowBRInZOVW3y6e4EflC8Y9v2S9L+NaX6vIwLw91a89rV2Tu2oORHfWZJVLuFPpNb
GdhsIKt2YDAua6T4l5YlOdtZQVP90J3Sg+i3k2+fY0Kg3Xoqt2sIoshcf650+gCYY4cNDWlsmghn
YXgq1racyyOaKiVrVR3Ceylze+IOD0om+t+0gcX0+vOTxHDhtn1LwmwMeYx6DpI+kTKpb+VKTeYs
NWtybtDo21ibId33IVIIr+CVOd62EibtNUKSZ83++F3HYL55KOgyRzePfa3agPWN2qO9bfdugXhm
+iFTs6JXw1MzAx5Fy64ZduGDk1FV79DtRXdRLEkEq9meSI43yE6Br8+NGOLISoxrZEwejHR6jsHj
M2cBVGoRl8INcwva8FDVIzmRfRND3uDFk2JZURCM4OxDfl8DO9bDIjrf90+tu1O8uiiIIkedCRcq
eauRPvWdSIfPgGZ4vUYvWNCT4JNHJVIC0wgiUxLfZ91kRLSNNVq97pL3RUCmQLdArtBmArzy2Jdg
E7paq2AQ6QPwTRm5gVDM0/wRSP9nsUzKIr+KDnMPNAODxTtUArmgPS/5Wn/rJGNBOirKVrwD6Aw/
J7eQi4Vyp+bWeo3IGu84gyfKHVGM/m/RDFMf6xzxoKegG7IkaghX8GCKm7mrg3JiMISU4M7N+OV+
nyRanlrZfCQk0FoWJ1v1PSs8MPbM678Pg+Ah8R6j6k5MShbEThVe5Qdpcz99n1Hmrxe/DusHz02s
VtoEEzLCKP45EuBexby+9bAoL9rAm+iBLzDy6sHxm0LqPjASRESzJkEbDzSChd3YNpBlR8ajJ0jz
sXyLjORDnmIyBgoXynQoxZ0pxmSF8rpmGhCBPEhEU3phu9JSJO7Pjw1CTDOr0qC2tjHHcuA0o/ZA
HBwAF5FSN+vNxFquM3mayCskfUV8eL9769MSMxXqCpf2zIOM4CEZF5kwdlB1qi4xdWzTeFXszUBL
EkE2PciHfbcsIo/aKHynjq3yWttiHHdONg9IFUU01Uz61KnSKFtDrL57Q5WIO7uB8SO7D62rpxQc
1FjOgBVuHrCB967OSlLToipLMmV3rSwIiH/7qMMnfh+BsULsUUZ3PjbEf2R6qLsiQLEf9QGfs+H9
8LVczAWylxZwdPtoVH/kW9fkz3fe3MX9xTZDSrqqHdPWJqYz4vt1h+TiEPDA8ze5emkrRGobIG9k
I88rjTBYRgA4gSIcy7fk607mN1EbIkAnPWSXCzBIm3uuYINv6HbL//A8pHrn07Jr/OirCdVcDmvM
1AVz52yJmWFVOWfV8ncb4k0oUZkVCtfeXkIpIkyFCBqEYlXGRRbMQXJSMg1Gd5aroqHk+z/cjaBc
5XgmNysKCHaMwlyFKX+1wl4iA+5+0yrCxCk/N9CWCjG/1xjhBQDVqPQkFCF9B1ZPCaO/t0Iacza7
H+4M+iKLtV/Vnb4bIkHhPDp60KFr80xYgxA5AhIIdLg9C1VeqnTJf0FgisZJTd5jAbJKtG2T+BHm
jY2Kf3hL8nIuQjBc+T1zT8iYJH5945SPPB2+ahgUGJ2Bkt50ReAzq65glXqMdXIf3S/IuYZoHO1M
d6ykB4dpnduEMkJdPfPJfsUSJpGECkYAxCMJNWwLxVVNUHcr615Th2DxiJ0npBE01JNvF3jQUkun
r+Hq15YYfrK/hBVt/C98ZpI/LLwVLOKoGwtAokLPZawJZobcmIGtclTLxg8bLxqodoFSWJMK8gdh
klSy5m4pdE4dDLXOVqAby4rC1c4ga0lev9Twh0p3MrQzu9c5AnueWgekpJlzgjZqzFgQV94WMpUd
MKuz0UrZFYuS34P5o/rWlXrhJMs6aKAvR9abGQViwkyREjOHNGE1mh4q+Cu325L0ZMpVsiEBUGXx
o15mijMxFnir505QyDy4ulzC+BF4v9E1GIP8VThflhEdNfv4LmgQnfffO87QIjm3MdGzbwYlCkYy
EODjP5z3QPeDVtCnXoExLwJZigLaojHmHF/n8qqt5NWHrVWz3Q1Ua+WcFMWk1KceGENq1q7Z5n0W
DDNFIG9W/gHFhpT9y/bGBqj+NTo4SWRew9IFNv99KSu+MSilwhyxH3E8fDA3AsP9KKSdK7yXiCR9
T6rjlJZeG0dd4SC5mzERiuGCPB4ZbM66mwU4aF1Ldy/xkuRCQMTZtUGCp7XqkbKJYqUxqV+hQIGA
zTOW1YeyBgz+wLdTq7MIKZe3moH9N3lOThWBrzTBt5ZfHLeiJcJ5R1/BCQ8ZkUqTS9dtfwlmGAGa
KojhZGaDB5WC0uKGMp0of4e+ZPrrM3OHr4Z90KCZOhGQz9m/BGQr3jSx8UJnzYoXFc2UWpnq2fUe
969bVY0eShdBJ3lI8ZbqR3i+V+pFXt3NuLpvC02xujPW65RyTjhhhD+K47FRN4Yq3uvz8CJh19WQ
99HQf0MyxMfWC+giwZd4e00qmjQLz4+rsUZzaAb8jrz8nMc3Bx2KzbetJvVPdrFSDb3U5RSkmVIz
KkfCU6U83dQSp34C44RqBmJ/1sLLRhxWYu5rRJEB/q7Pwe4cmFIvZXRavebV9ulsqKuVAg/JJM01
cQrDPOXwRwGA5yJy+IhuAQQh0Gxst6N77gsLyOa3JEU3xrM1s9E19q9TpVrZidZmSuivP1NbhrTY
x5BaEeWyUOdj1+HkiyOCUv1tVm0d5AtpYoih10CLnPDV96tWwcipas+CGqcF7Czi3Nu0s1QFiC4J
pqMM5hvxqAFn8KvpfJNgy0cxmE8BHJBi7gm9C1S8uEkUBEUaDEeT1m7kq2KAIuNLQpcj0Evrqikb
f35qkMrOcE9abIGq4hV/UW9gOBj8LYTIyJeDed9S6Q0LmHmueUgcO+8YiOHYx8NUNT+NqFdRWGr8
l7zxomeHJT9/uGqXql++B4fK9U1gbL4AuPGbYuCe/Fe22cUptxE4ARKlaRTP1pWaovtStzKo1pC7
WZhQrCmjqlWdhVw29tgaSSI47m9HC+uCq36uyHIBdbPVzcKl0rxiIVvTWbUUD/wpgkKxZgTg1SkL
5KZzaFtwGTvqpUaVcqLzcvj3WWl9o+mBm7rDBAFuMUrgq/oqb0iy0Kc8srrHQIZ0Qo8OglOmtPIw
c/qAKAGZG4TkQsR4cPoOqVlcFKJuM8nk5jXlI+GmAgTkdnW4N5ayAahbBD/Iv5LDOT1W6109qeB+
3X8vD7fW9DqS1FE75F0rOdS0WELB1tHmWlXCrCSBb7g2HGdH88fzSZ2uG8ttHTrDKts54LruspG2
vTD43uNSiuLGhBXc2DgSpQsniwuuGTvY+Np2er34UgwdNXKqBHPmlRqorAtgj+XdpgbsYZH7vtoj
knsRU02gNgiO8QmCcls3MNwlIT0i1FNe62jncZHxdvd9CA8DBzOv0JghkDEus0cxsBsumNom1Kp/
e4BCKkv93ZEsfK0+cIpZ1Trghua09IgyM5DEKRUWTspbuusjfj0R+K6HifH6mE0BAXChMyBepUjE
7TzuZUA/BOkwyHwFUeh3ec2jpCwAYegQt9ktWJyFoFNpWtvooYbJspZlI3AAIPrvsV1K33b+q8BI
HDLtmussTpArQQmWOyqrA+EZgCFS7rVNdMCfrNlrfvcnw9O/j6nGngZngj6XlX4P6Iqz8AQ5ly7Y
Div5TedbHEanE/fQC4QyNHagGfTl9cXsARu+A8XLP1b1ymAjsDQTdouz99rXwM++0NXnhKrT7GmL
BuimH0xNfbY6zdS01Msu2BzzD/6T1ilfI6bti0wogT4dbtp3Y4hu4+3DnWkL85hWmNojqwO3C5Y5
cYOPldaQnhJeE6X7bjGdJTZf+juEnKJBCS4St9yeUU5T+iv/zrlBZDkOUUN9HFyd7xydZd8ojQS+
EaKk6+0T7+Eg07i/31FWOf7vNklhc6BTt9qsUoK3kcOBYZr0rtECOL7bgiCC8Fgi83QeXH3H13Cb
cq8qB7Ur7xRBlxA11HpJVO/10jKgGYf6WluN9BRNTRaNcHVUfVuEJNYplbZ0U9KVCwzhtCGyD3oI
if64SJ3ax/+7q71dK4RW2mUFKw3dJwHKR8mlptSgABEGVs8yJb+kazVpyp25SVHd+URItS9Qqanc
AXEwt1eFyGcYRERpCk9w/wn32eAqAp97rOLx1761rU4wIIXxTCJWHX6aUVnAHWokTCdZyOtnyWNA
Psn8R2A+eFA/o1JzEPvmzYyWs3dmJSPmPckS8ckhDUcKp4R1hmfFCn/PSgZTAPkHows32lN9hdte
wu3uCoTnwFTIe3g+UV1QTF7uqjiH1JgNeHxfUAjHS4wEhumck4wHiinTv3GXWwbZUclEJn36j/fe
bh8wWlj4mdd9T2b48S/803zuYhEHaGoCb0teSVyzRtKkVVZLsTXD8NC/GMwUysJpQl3OMfRY/9//
cg5Fv6qb8QthI6hg7fVYx98+KaezRD4lR1Whxo+hjwNuag5CYSOmPB7vJl2KFMCIasY/dkU4uwwX
OgOxmZPSiYHsBdBjQo8WLX6AB3B/FkrX5kKdKRYlfGuN+LSmUo2rPrDzZvMAkDJPE2+tFH+j86KG
GIBRGKzz2cHpzttyCCbNP5QfmV8IY6f/1ZA9vCJMFRNjkBYYmArwHyx7esvc85KfKGiilPzc+iYh
+/uxdkq/Q9C0xBLeHvmLyl52BYo+U0KYTiUhZDJSljA8wGWkl0KeMJb+CptC21fJ9u0FbCfS815g
F4KfLk+KmmRklLpNYughmj9oT8ZfoTalrtTOfxxSRIxZI11hApRRca6mD4xJ/yR459uz769hFOKA
pu9zaZqvxiXgvWc3GwWrYN8KUbWfLLZibaNMiS7VodpYtkjjqFfPYoeijAQEk5/+rCQMIWbq5Rqv
etYvSUKU41DIHKf4rE00B1jnIUEZ0kGa9OBqcKUlarj72748axIFwMKF5cI55w8feGuxvv9RISbb
m3j5ag9WJ+vzrBYyHi2XP+uffUxzqgzcvyHOJ5pWYKCqRLXIKWTv4TNaXzWmSKxJMzQdahPI7wxF
6ZS80vMe0MdWgriVcSBBO8LLon1g79o8TRXOD6Gkkv62WKZ5VuWkzHT4a7WPusuPrqXDBiud+wTV
6Ha8KUntjz6KCt6U+vdZWWqiCxHY+BEN4J0E545aaB2Ic7t33LXzqyrQUJ+XzsxC2qZrRkA2aR26
n7ARZs8IlxgzUGSUwRssub5cK9A97xnZZP27TBGQB/DZtEm+rxMcfQFVyPuPkaPyaNoNsOswbafz
Rt6YlhinR8bzZtOvEMtEk/fIELTRQijLWINheavOel19qBZWHU7BnILrQ58gZRiSrQijmHEb+NxG
6uDjJD+4FNfxJhOdV8bhFuodmKnRbffMZl22HzD59AlMaFDdS4H10t6Cu/DHd4LaC5ATPEsDKFNy
cmQdli43FADQ56RP6KBja8ln09zmaNrkpwjQnxXG5M0SXihfTAsQAt84G90jdqSnmTXVdBbOj76N
8SYk3f1i4Id/Ox0ab5t5c9H/FcFy4GExlxgoa+KLqd+W9w3QMngvWE+u7zyHsmO+fdYz9f+1mlEP
UuPKIxSBhkYzsBfX47RzYE84dguG1QeObksTsM4JbvADxLAOfcFHG20JgKEceBDQsudTqQ+2hYSL
EvOKNfS8uGRQ5pN6lbmSUQEMdskSbLFIceRwHfK7LTSdhU/0Xy+omAeu9jfGvd2Y+1Iee6vAnE5K
tn+roFZNca91iloohJK60ZJu1RlG4uanBHabDsYDoai7Z7vptUPQDgVRSJERr3x9PhOdYVtmX983
WJmj7qQ9FqTpsnnGSXQVMr2NZb3lb6ohtfO7oun1qqyBWLL95App5vM90QqHfVdmyipGF6cRerhL
0YVtrmn7gzwWSThrTN4hPQeVUABuOcJ3LkcMklPBQgeasz/DfFSXeYyTfjBRHBVtneR6ipWPxoNy
RuNQ9tT4gc6WPaZva1soZNSlJueD7GEh0InTfsjfzcsFsh41jtq5TsZuJdzVCVR7nMfbCM6M1be3
eTYoT9NHPCYhaR/Tg4bJqShb2VMLNt4YIR5aBR8LumKrIYA8j/gUntsEKqSNNGQv1oMXODhLjyX9
OoNrXXBNxGuVXi9r1rVaw9UCP3t1OyhYzWAG/6RoRkw/CIqAuwdQbfgAsn4+vsvbal9RMoyeYg3C
SL9x0AvUnYttfaSjwVm4T8FxllE2XeKENd5rSuNbVm9/2mnnx7FlV+eqz+a5fWod+u344Rk7xKWX
q+vhBoztJKDqhyTyUChVcUCV4V30VphVWDwelCpHmTeHsSC5rAThEVi/Ff9aUNQqMdw4fjVKlL4l
ah5fESlJpHk15UffzxDY73ZnMBS3RMsDyJc6KqJCeTK7wf+KSrUUAMP5i8YY6D+QmLaI8ggJD4Cv
Pi+29IUIDHYaDjM7sSTlcGxEwsRwLM77dBuxb7Ggm4TlTuHqZqrYWc9e2/Dqx+DbLPKk0xvnWzKF
lOl0wOLhLh63esF7wg8Eea+oIl2rTSDENCBRAon65QLcLBoji1i/x/EBibP5Ly2tZTHFbJqIf2PN
w33s91Vc5DXYo8tJm41f+FUC1mpFxKI3yZWpLYmgzSqOuhA4WexXQQpXg8OGzxKu3vUffozrYelK
CM2ft30G1lvIFgyeonadMgj0oUmsBa+UW476i/b/g0E76l8sEfDBEhM+zssWRxBXn/Q4GGT9o6eC
BnEeCe4MTMUOeMDON6wwW82VyTFBfz9BMrygf/0tGCiaLO8ZKYmw+sewz8YBkjl14TI6eOn07uaw
h4hrEb2dF/wABRVF4D1I9G0uwO7GHYMZ092O19UYFFJjapoweCGoXF0kb8n/m5I8g1B+uVz7chnc
6r8LGA5qWoCV4gu0MBPEImUlUSyHyzGUfKAt5ERpkEpymn2+IZY+dtxh+3cC9DK8jKv5/ic9Q0+R
9meY8pGMkoRLhsXF5Q5F2hO7q7sjvocBpadhIz03TS4jUWvFf/DTOJGJsGOfvlf1oNLRGgnjBOAZ
Za6pkE4DrOOG8xmy7b4l51vD4AdkXeXTkWtuLEtyWOGoWomG/lFyjx7r3lmIiW5CmX6m0B+Ukl7w
LS6RuJ8nO55mxtwx7aPjdQXy5Q0QGZuV5D8axNv+tDNj6wOZG3Be32NfuRu9Gqt2Bf6Z9JrPQBnS
X1gn6MLO5qp+MSjvVFS70vzilWMRNY28qtaSxst8ZkM8sqzSEhpVJv3ixX9wXE5MrnxxgYOxNQ8R
4APIuEoABSRXlUR34Xy1J3JfJpmJJPgAdFfygSCtpafakpVmIdyKyxgXCCQ72F7TdCG0Zc9dHmTL
oqu0LpZmMa0TaFM9U0TdyWUuhsgVJAwzW1t8cUGCa1bq789lCWSQiy32UN6HQjFHMRdlN7gKshOo
kGAmAM2hgveGRfX2W2wmbuYxqhO0ktBTkQmiJek+oXjuMablb5A572Qik2Vs/5rSjPtHDgoKg0YT
CKwPYC1YWZn8GPMQ1qCdQSx+v061yNixWl/+1rzIA32gx8gPmDAWb5vAoaJInw8wX1FD+R43jt0x
JkGULPz/zQ3g4HQsrGz8b/UpIB/v1tGBli8amr/u+//ahxolKQiOM1kn4LjLLEnc1mWN3c2Fv1Bi
qMWk8xdDzIuFlIHq9efKgequVYPl57f0+Vb9LpUXO3dy7oVRffeTyzG3e9lzlGScG1uG3tf8YWbT
606kU77gaIbwhRbe8wszDhayniIbe1ftVaFg1byHr0KhVa++11e7U8MTwFo0di2IaW3/hYFfxlRU
J4nhI4MrFEi1D2uL3YKVturxA9QrqNSB05rz3CF5qy6qyLN64KJ6bOv2UBCwXXgCNZ0uQVEb8jUe
tD0XTsZwQ7vDUPnoeF1fKrE+Hz+NUrgxmvPwqhwFX6hbGZcpzqM+iBQRmR3YfAiY0xESpRJ5FiOX
C0Ez0ZO6ZOVvlcQXdPmZWn1wiVqiMXiPIGCefgDHkVEGPKSnz+SsqoT+OP2HhhKbFRrv7UVNX7W6
Gyp6Xd6wJ2ZwSrArkzNO9Wbc49ii4nIPt5fNUys7XsI2lR4lvVpNGU7XjleQW4JnYeazLxSILjy3
ryviyIFUrQMmzG8uwmx/x3QrDTt1WHb4LhZ+L5DQCuGJYXTvyX64EqgmlVuBsMciPe1fZeCz1HRh
MCqXrAr6gXOgwtB3ZE11cxiCDDJ0ogS7J1UWpx11/my7fi+2W0BSQiVVqQwgSalyPTXyE46DF0cK
bX5aYvB6E20zIye8YAgzghW28ZJiOoVHb29dNA9ehppGh/1Oaxp/BubDpogAIS3j6Z5Vq7NM/tK3
c8EGKjEShezd+eb4WuX/bFpQi8Tv7Fgd1aJ60PaqTB/4MrYTVMBTKZqGZl8J+NOY1zw2WFT6zY6s
w2xV/tJDYOqFtGV2xDvGIxQBaw/n+7Cy1+P5rPEMBoKXm/+HBf3YqGuWJ/UyQxbI/vumHeqSKOuN
iCx9U+2ma0XRvdl041A4xmfCEmedc6cD4B2s2ao7ziQxL9xAhjtwJBg1F1PGL/tuSs4JO+V3hEll
L+LXJp2R2Pkutr6aBWY20IAmjGMIv4gMqtGhtHKRKRMPrIKJXybEU1y89UoSWV5Ga9YlsIwd5rRz
EtofWK6ehxI7ZBqUZzfCmv616keUEKkE357hQB31OIMlWAf3fDWD9ddwCgVrQcthFmrzKa8eDGL0
qiNF0HCqPkgkyTs6sUXu2dEJjveR3xEv5Zq8QtbV3cxAlSFKhIvb+OOCkBzcSJ7NhiICrnH0HQZ5
2VK9kNtlJNJa4WaADJdGKVsm/SnYaKwtrkCf4aTOqFmIgBxi0E6SrNoQxcVhTZcx3eDyTV5FFzlj
ktGoidI3oQYdgtdkDXpawKBWGtqUEOWi5n29aODIyxnjIwyIRSQCMvR51E0XhyfEVeR20xtLrVu+
9L4MQegHT9E21QEfSuOXH6r073xYgZwEnHCcUo6vdW3WAcXXsKzQHpq4z4RWzHYjTDmFux2T5xX1
LpnnbemPu4hVFY9pxKRG6mtyZjkm8F0BLMBy2D/qIyfyQkVb5POfuwESdqgIhllVlTNpGU1uVzU6
6QkSwqwhPZbRXAeq8fK6jhRKjXupHXMFKsFvvPtVlG+EAs5mEa54g5jFrnJDBdpRU/l0VFfGWHdN
qypaaOwkAUGjbR/EHDIDaiXjhQqxECkZrcm+gicRdZcLdM6yjo2F9sK4rTz0tCycCGxaQ8AJEcee
16a08b3X0Ocb3zc9mh0pgLUrFUR5wFgFxlKj/7bzJl0LdBRTe9kd4vn2vvYGlr1ZQgRuR+CLwVpP
8yy/Q2al2M/HSMVe+5Qws7CUFMHBy+LoO8YCryikIlRj9bVhQ9t7IpPBT8+/8qs9TxgU+AnZd9yM
5R3Nxm8HU0HxJelLItqJ/+0IO6Z46ZKaSuqZ2xRq6Y4YWY8GTTTcNzkpFsKaZ0X5ZvRQUkgUOOG4
uLhHRJOkW42gQSSVY+Sp+a+UcfdRx6pDKZ4DeD+Od0RThq2IC2uK69nbcZ+Jjd/X2QOZUOs3E+SQ
XtpcQJhS0TyCipLghj3ZVchnU7ZgwlURjqMXiir5M/wCX2/sI8uaniVVuSYupx2r10XwD8OuSRIg
v2qcNG8xvU9JeBoPGtHYVwEDU3E59h9jd/Oc6kYCRdxa8Lw8jl7xej4VvWESvgB6aSnbpGaZwOD0
uaJl8yQXcJeb4T4s/7grBi0w+1rpMd7uKt6QiF2OH7WO8A5bdR3+NLKTFz3O1nb930q5KokiShqw
CNWtyJENJmYaV+gQX+VGrmn8zKE/PV0K/b6dQVKnYOB26pw53GguiZ3jo5GM5Xq+6Zl2Rc6ZGgAh
Ux3bN8OuqcmcDPAXNTkcTu/I3e5x9K8fCialmAOvxduhYPZSNzhoesb+GLgBQ0YdY4kWB2FBXjsq
aFb/u5lLsAYqIHgQ8F/VC6rtTRwg+h1noNIfURlxezrs5170ZISTPz5xmZ7PJxa9GWLUZ9gacCMU
WMixxqXBDJo7AVl/3cVOldZmmKFg54B4izOgc96ZYj1/N6nyabOLrMDl3/nrdZcM+pXoV/0pQ4G7
hCyiWN97MgE7WF5DpBj4Et6NcYbNOtZJmTDrfChmWDEnzboayRUp5rI4+xFotvQKH3XhljOih8gP
Owz5xaqv+Zj1SnzcGBkgYNEX9ww5VwlXRrUzuCoa4AOgz6kjG57yJhggnjjNS6G4s4aulFI4gDaU
Yw/PwGawO2o4RdJJqcGO1hBW0zPtLuplH+EItNZMm58wgv+UWVpGvqI4zJEKXuVe2qP4tt8uzQow
tNmDJrjUIbmd420qsGh8MufbwWnRLhKDu72iT/YxgCkDsoYLyWVYGMdoU+t+A///d9f8Gcjhw+IV
O9Vpttt6XFgL0mfYrkhRGB+eS4zdMSSI/Yr5JEe1ClCLnx8dlHdhqffBKoUYklbT8mMJoPnMOkLD
kQIJYbDF4eTux7HPL5yoihW7keka6NGYu4xeK+R1qMCEG2K/lWDDYWMUu/5Sjcnk83WTWzIJWFiU
6oCPDVfkYAzMTxZhoLWEGPy9bhVBjeBkZQ/W5pwyHirLecC9PlKhlPLIqvWU+QxJDTmNa8AppCsp
Hr3vaNrjASpsTSRFQ/TQhVGs4DvQlGEuitPcClczhDOqQupUiwKUZ/uaGeGMAh5WvGV0aZBfTduq
77aWqhexgNJe9VBFUZBh4/o7HFTho4az8+ZAIkusWzg45hmqOrYqGfN+eGIdTydnQVyOYXcVzNYN
Ft9Jcnv/yQMCV1cE0sKY23FVGWlwGBhfjpL347WowG5viF6MMaj9D+WlTeWZRUS7R7B+KkbYEO/t
WNoTKmJO3NWf83tgvuUe3lt83LS1+pNcx3g4fdgXBznslC4GfhmRqXRVPbVOqf6d6hsDJSBg7e/g
BGrYo/ak5LQYj9c9cWza7FfTUEGM9HFK6WNhmG5/ZVKIzgfkaYOEdPtv+LIjKLWe/dzWkDYJhW+a
XIcV+YYuYxn+jGidZr6ibifZT52ahyg17WX64dubbGpq7PxRTAlb4tfrumzBFugsXFJdpkfqwdrs
m38vKRFh10iucWkDHMiFhfWeIkQ0w54V6prUzTYdjRH8HGdInzHctVDpkLeajb/Fm+QaAzTRCz8m
ZTmNIR78MUoLO2bKBW41fzQTSFhJma4V8NZufwoxA25GFO+Nvk0sbEpd3AZ4OffeJb39ec370NaW
OLJolDW1R79FFUZJGDFPtepd8WC3tFwZxFYXJVcOx/UsLt3457uCA4fDWQJR2LPBqmimzEv6qN0N
bMN32msvYR1a6q+BnxQ/taMGfeVz3rcyZJs0kgrmSG1nYR9DBIdLIY+egydJ9/qmYfRDKrRamo9p
nsOJaPFvH3zCI5Xt70NOSG3YuWvgpjAyJMrm0AMKRY4KAivUa876A/Zb+bLPqRM1EJw6Rt1vOFKi
ONVTWLcHHK6dxgKywknmtcWu6XNWBiUO+9GaybCddKjzsZJ4N8MT1yjJMaFtGZxN9CnKE8+XBpXz
7U6vXvH4SA1WuCh0c1cdcgUeQwv9uqsP7PZNlKLBIFQahNzwa7cAZ9EDgTr+vmwsHDThm2vV8CGm
93zRxzMPm9r3KwRsUNm3r1Bbd0MzUyxbYF4nK6VEec2VR84TTri5GRuyOeLyFQTnud223lxv6JnG
6IHPzNHMihI82bFUlRt2t6w2Cm9OK2yskYFQagp6W6k0YSplWnzuYUKXZ2+Xe9ZY6rbZ/eaFgGrX
xM5kUlYtuWdktNtKubbbtZHoVeiVrunTGeLoun1uNX/Bf5h8W12r8AuQm4H9uBnZg4a6Vn1C5Yjw
rTvs9woFGUjUPvXyg5Q75PFR8Jf+X00dmC22VTWL5xUey+DUNI/xJsGSZ2dNq1UN4AArsOv026Q3
yCN37tMZC68grU0z2oAovRUg8AY4GElqpM7+zdffdQUJ0/1ylkfju33NFqvOgcPLcNCdqvvY9/gf
wrueWViW5TgDkMWiFVejhnbfNbwVvSekLVvPrvEmFqKDwBfONGYEkoAbYDlcd7IbW69+kFeV4Y3P
lh6oXF2oQ1VQIoYXaOR7RCUloOBdVkSxv2KlREygLtvPTcwO9WkBWm7p9t3pvFfMc7TWpoHrWvr7
OmOYe5ihFRHwDbowPL+m0oEfvxHcH5voLn+CmtFsin7p6riLGzQn25i7320NUZQCjhaiRVR9G3Z5
S7T3ZwVWycVyB30f63bVl0Fl3daxI6LBCq0SoagZOPHFCQCYd15MPVAy53sfEDN6vtRsrYUdI42G
jvOFI8tZJL97CuKTQYA7HV688Zr+QiCdWlxXvQOTPSOrpaFxwODIGuxSkO2I4hQeZpYlybPMGLWD
yAoR73DRzoRN4ApqkZCh4DnL9ys8NiAUnY1QLcS5gT5j0QTQMAipohmLmOFm6dQzqJblj0HgtvTJ
fX1dwici3HwO5IBK6P9ucVNut6KuOc1xg7I8v1/rKKQuKo3e4aJi4r8/TVHsSq0/UWLCCa0HGvAu
tYxPkxb1EcDo699bNpQ0nlqrzZipGH6upRyyR/VRVYHZa9GcOsL0h6gxok5ebipG3IztFta0qioT
OlUb73g4Qzf7U+yfPobWpgu+prROT0EhJGvM/+afzZvbishMOfJxF9WPTF2vFHXTXz+cyKW07nLQ
jfSn4t3H0fbWrStoJC9dtAy4GCXEXkaBqjJRSKi8cDEfg4swV780fOg7sIdT+v9kkF6VjMo0nTJq
kJQ49dt2lKiJZ37g6PKSFBfciakVhG7AHgDNCJ80n069RcUSlcs4UnwR3EInOctHEQ5wDhbEHSDj
kQYfRz/MCb9c5h03RMZfb8OxVPS76Lg0yVTqzTE+5ADHWH8Ww6BP/pwZhAww/KpLsAz9m1fK3zdC
P/H5LqeuVQy3DPXx1EvqKrVZGNBgr4tl9kHrjuY9sZq8Ru9SqbYf9Aptna5pnR0Odo+P14oQGiYp
q3qPZ0ZQV+7KjBFRiTIjrbQWww+Enfav7qLpT/GX/WOTSBwsxgNh62H7QpfQWUcM0ASoxjsg9I1c
k4qSwFwuZXMFRZJ/izMskThOkedZ4fe+8Rr7BrM/lxwlZAwrT4Cn10djNHKQoFk5gAZcdN+xmCpV
0RdVSTpHuH03vAIKOLoLB6mzdXRKuYoDU6yJos5wS+wzRkIq0PnxwyKL5FUP7t8vSXdQ4zTLPboT
HSA/OCa11NSjEOszMT4FExUcXd8O9KL50xLadZ4Ys4rGlI10iKUVNP/s/0Yk3GEcGVW2S6PyobjL
mVr9LztJ7ephvE2T3SIweYjdNk8bXRMwORdQr+VVz/u17aonKUEVMClqfilPplGsXlVkGcEhmgkG
FKKEe1O47uCALkpuT8OIwHpxyZ9jzE4I2ygXBye9eBTL1HdMjoGtKragHC9EeUmMtC/18Lj/zgka
n3XdF1oxuepZ/DFqaeQXfj+GifU0j0n1eN62+Pw6Fb06krD7ZxIZpIBro+h/L1+nDxibucRiU8es
3tkQL4QzMfAgSUOFvosTm0IbmrELsu3SWe2u3WWOrAv1WcyFcKFeBwEC0QjAHGTqx2oZEZ4JxukF
b1vZH5SgVpDn1A8aHp/+tQj+MYa9bidpYKhFGatD+vHg7qQ7ljW93xyVRtn4gId89QLJdsVvQ8rq
LNs/k49TNFHpIy5UbqoDySbgTvulKRMHN4ryFcMjRxGPpLuUnJIdG+w0dOl0Afff8dRtmfcNbw9G
ClB/Up789ajapofv2X67uXkVNOMei0J9v9mmI3RsG/t2A1VNFHaZ/O/WMPO1Woj0bW4mFLpWSmMX
aHCaRzvc48/v0hTOqNrnbksgIhtG/e5EwaynSRC6aW6TOx2Bve5dGbocq15unSbuySlKCTZMfYYS
lhoTjslfw5ytkmOSlAyCwBUK4VbotGSMCcXfmfiGQ6TlXhOOUEbCNyNRaadSm8kPNBkeHGqQGGYB
0tBq9awsh/mivU0lYCod5VDEDNcV49z/9Ue5T9ejMWM6yCnNQnWoCZqp8bHtpO2Fa6nAmpUEw6Hj
Hd4T4BKF6KOkDu1sI2W/z0cSUWvf50bLfOkmykOSONrc1wbiMgtQJ5NBTlV1SjmyiQwC0oWIT359
WHeq0z2V6/gxAX/MeIFYUOYSFGC7T6eAGigatsgRBJpIr1a3XsKRH3ocvqReLMBANK2xTBMVMMMv
zpKnKJnJXGs9bLtST4l7ZorRMQFrHIS52yCUO6CMG7hBEdEIUq8JkmtxLTLk3JJlwBaT8JzplJpH
1eGDIDD4/2k5C5Ea2SB70dTODhFr3ljax0kAYIgmZqnDxTRNUdjZjYk6T9qVZZAEjuLKCib3WuKC
gfbu2CXFrdLEKXDzup1YhD2+Ib0wAZbIizlJmusIQltVmKTT8p8PaJjbLLzc/OIOaeZRNsBRPrP6
8PvzWQXCQmZTYJhJVXdi2t2yPfmL+niqZAbWx3bvtH3H2PXhMqCnwbQBKxI2UsJ8ADTLMKmB4UXn
9uqvIsp0aH9jSyc6DDpjJt8bfsmP5Hbf5B5chWASq1BNlEz6vhkP3eXmIJKUTiYqfimVcZ3iaH3i
9OAM1qwSn3IJDmPp0xR0I/eNi8nLa30RwvFlyWtcvLXjFLRo0/t9wrkxo2WFT0IXQD5gs8a5wkfX
94C8U6D4v6S2kNBKh6KrNRJov/Exey/SsR5gWGvYSoWctCJchkDq3U2fc42H6reBglS2d7pUwocS
y1KIwdzNJ0/0W/irjLUJIR/EPSTMpEZL7Xf/Juj7rMyZUULn/Laqfv8X88rFng9B9G5YnoAVtHls
+pCtsOdmNiyOm1plgNVcOWIXhQ0rgS9jljf33hE8hU8cSnS5YaA44kU90KcHs6T3WTs+26z3am+2
NTQaH2TFjoap1kA/nG8extOQmNs/dqpugdi61jHpARgCTYFjKGpJraICp9jMib+Y590pj4kv9DWV
coYtGOfuC8EoEFPHNkojnBfcjV2U0qHYJPlDtBBLNwWhBHnXPTeamgSfELRij39Uqpp7Kw3q9arQ
A/0Z8uVVisA4DZWsUiF7pfgDGO5O7ssfdXzLDqvk8t03a/Tn7/37e8Vnlgz+WIxFl0DmyKs75juM
Y0ZGLD6Ft50BlOID9+fI2MUG1DDyj1d2oz3O9VSvvcvaNhtDuuOUr++WNMN5narPCs2laAmxa15O
FSZilfSbdkhIYW07/xY7Xfq3uizDFzsuZfA7I8jztJ453FpNxEoA9R192WC/D23G+GXF1IpGEp0f
nwZh2JjuMlZYImckGUIsENQR/1W9hJp5buFB1rVhwFbBvPIeZjlzugUcAQKd4FYUaCP8v29dZKMV
RkEHIbnNZA40Hh/y/xztRl9rtmbEfU8MkFPze9t4XCZlhKYGW39/Q30dlnrmKPJa+QxhRJaA1YPg
07kMf0a10eIJ+PGei1M1Cvu6FVatIXYPDaUPv6njOCZlBnIYzjxOByxxXG+SOFD3poQoy8nkRzJx
NfrLxHK+QmZ+Y1+iqRNd0CR2RAx2Bvp9eL8Rl+33uCkqv0KtquMTqKnu90ovvS5+LLyUOJx74QXy
EIRaCUvv3Fx2uULPbzS56pYJyv6cqkLASUhBAjf8hJc9lN4OXASjWr8I4nx4MJrwXPBoGcMZMD5p
oeNdCQZT7dUrmf4N5oxrhiMHh+rqEtWtstB72nalxnm1M7+bI5jlsjNJm0RGxsTWg8AQUQ7nJ4x5
zKNOzbZKUS6iBoeUpxqmgr8sULeFyeJZfByQfH8G/OnMv5XnWsl31uvI3sCZgWFS3pH/y1YRmAs9
LzB9iHlv7CYEPJAf+jLJOPirOsePStvmPUjWo/DeoIpBlzqoQcrgqYbVKIClQ0IbCkeiJT1N6kpa
R+Ie2BrQDkOsSZzfHp9aiDR4yFrT3WNkLqqXfcdKhVHtIb3IocyEltvqeaRRr6E3tEAWI2ngwIEv
Q+IirNOQv39OC58pbVd1jP/vr4nXWrkhSxmCZfnL3xA3ySmWe1H0oSmmc2ptXUdqKHneCbzZHQYn
sXA8C7fMPIRrT2Ht/FMt9GNsMsc0Vag9VFAMUbFEfAb1azTa6/hXmXYCtTZOgx00gmC3epj2/yVx
aO6Lm5jlJW5s8TIwIp3l+MoBWYj1f8eOE/rScxt+vCS9WGfcUz5qT61iBrwPTdXgwnb3f5/LKM1j
Y5gR7UYTtb6D6xHXdGgh+2/GrPd0Q6lSWsCarZM/YVUxa8lmVu9y14sNQWMdBSiy/D7UcfX0Lu+J
EbubMA3/SUClTle4GRf9LwTy5wZwEx4kh89MipikCstvsn5OI3Nwze3k/1v2zseUsKvr8avAAUxd
rPZHlY7NiyMXWsrKkyPQJZDCA0v0A8nvtRwAShT8+komMpk6dRg0JipCuR6g97i2NZ8/0zUWwvkW
HGd/CieDJ+rJ2WitRI8A7gU6ptKRK7RvgiXxRsfi3wAmkiASrXqIYNHZBJOqEJMLvJ3HgvokPt8w
dTN9ZK2hf4GTrP5KSExWX1QGdXKFbsUOcUcYGj2robKW3Jy97E9T1YcSAYHmnspEFGCZhaB2ZCp4
lu/CcsCXMaxGdgtjBPzkEBv/sKeuCoEihwzbOAW9dN7xSdpSN/T9szqM8kJRDXVSvTuwhY7dCRf1
5XKQHlVMA1/4Sc1mMVV7yjnCX75unRso1+wrUOs3mm4XtszIfiual4xnDIE3U6DOm2hM0RUh9pSz
KoONyiQk0lx0s1BgQUgqpWyozzvT8BP9ZEnaSQ8qe0d3Qz1XbCPeZnR3uWvW5ppe0f/SWLPasRZm
DqLZXiwfeHPqKHy0+EUDog9asr1lcVi3LgcqRbT66WNtN7Jom10m684qISX2VPtWcT+XsK8C+TML
O0G2YgT7DDTAL5T4NlWHQgtksSkhMlSwGChW/WMOUhJlXj5DdKMzcoTLFdD20oxyY/eB9nU6Zbbb
zIJ9xC5Vg/pf/AzqbgSFAImpiNmr4g+rcFG2dH7KaEvMhhZysMsp2Ujs2bQRvY1jOuGOehqvaLZi
ttWW1ox9l2iO2vfACb91hbLJW3RAijEjgBCCFsMooGCtJxPlX9PcmvsshYfnnuRQc2PRIgKXDPHu
7cMWQBcxN3Df1+QNmz04pjWlloC9sy966dv8m5P1yMuIl4iBMYuLoiPOtoxJO/rW2vMM/W36sAqk
ee+PnR05vDmzIh14YMAhM+87A/LccqcquJnbg+3XiJFjf7G8glkgr34ApUBfSU2mmmaw6LTcadUN
hQsgoDFpPv9mz28JZKSTGmvX8WUzPkycpruK3IaryjPjCV3B92TdaUWJxK/QQkdok/e4QU13YjxN
Gi4HIZo7qu7mOu9ti2Rb81YPqjozHJWVy6rccYYlIlRraT52seILmwouKBLuY/3cI7J8HVZCM72k
xR40oOhg3GEbcPVjd7+KQMDVgDR4YhBiMoUgksCFV8fyYIT/3JG8Aa3xC6EnOvHVRVlnnzmVoIl7
dXol/1DMatC31fVmLRJLlNQxNGrjKY3DImGm9WRA0KHhI7z1uvllg9EFb+yCin9h24rg3tQlw9lU
gFstQ06/pDfOS/QcVADFKrReE9bSZaSTwMjh305U61QVVrSagDI9Quzf8lUOtydBG+nmGumRvV9B
4/jb84KZLHDwSrY5tR4roNXkTcte9T4aY2W8eWofeLkkFDaHDWvwy+3EsZr0ecuFb1hlpfrXxhBH
5EwYzsVhbfa29lNstbY7+NuwwF1uKAQ5joL90II3Avwe9feUWKKwoMzxhgg0hkqs9KYctj3ze5f1
hEdxkwzrlpo43o3PZtUHED1c0UqZeUY6NPPC3iZYzkbx6wRcKfEgmd2i8QDTf1VmQbCVrHACj9F5
2QbaEVtmsLJXnwL3Aa0ALD21BPj2/3qHqIfjmUzYJ7XQtS6+yAR1hGnEsQPNuozL2RxgaCh13fcp
CacpQYdhwqeR7hihv4pEqGeORmcdX0U588SnRL5fPeiWRsruhDKJuh9qEHnUHsBMzdt32ezyfDnD
EN7hi/O/E6R+0emHQrNXlQe6avOKvNiCYP3/NLO2zE9sJ6VxCy8dcJork6vHJ5MYb+0Zb0SOwyey
+rozvMEu3IGt4u9grvy/h9814pNH6nraRkSpuoTbE2f+XwjyElLNHFZp0CmOqk5rgAK0IHRznPZG
SkMLw3ujFG9fCpxyePZGKDX1eWW3nRfD/xAgAqtHxljw61a4VYxCOcqKFivHvsEHah82i+vM6JnR
X7dzvOjQRLrTN6OkKOKC87yDkyVEylmo8BxuWorp4WE1HmBYYaljXVup71qk7B1/ofFf+Md2lqkT
lG89RiYZEOG1U8sLgxSbtWYfF2NusVbzB4YnR5QGF/NZsGHINtG87pSnfId0quZw7ICeN1EUEC9T
Zc+khYkXBBduzFa1G/wm60P8M0PpNM+VSppKMlelJndRUno2oKxPlXUoEHIEnrSKsv9ZSwzdUWNZ
xQzODh6uPlPQOEXYj7DcNrFcyU7kcSztmF031aZlQ5/NERBnREwzPb4+AJAbwsKp5ycmuip6v+ls
DcswkRlh33o1eB61LnEl6UpxdPaWhRv9cIYMbhzmqKgjHMmig4viHQ/qshNOIdJ5RFBEU8PeOHeY
HQmE3fDcPcLsRzqv54d3WG84CcJD5ljVtTBXBceIY2NZrb6Qkgt490NA21iS04Vf+6CLTrUA2kwM
c/LZp3u9XwWz02Lpc8dSb6wXXpX9fU8TO5nQsgeW7csddLf5LJeuLgHKrrUJPw8+/dnzyh3a2Bo+
/4SSGB/M8gowwul/HjEqLLyrTO7fjlfEoY2uivxjZbNAD39flL5uu1ePBZtEiOQedz3H4KlSPbs6
f7d9kX1w5Z9mr2Q+wMKmpBDs9mlsbvUeaS6cTQ8JKMo+OfGLLUIz6c+2ouY4yH+RNH/+2jQIN1zE
TdPlQ6IXf2WwVcUKYj9DiFgFhD+w2w1s18ZWlvhhkq4qlABlBSp0f9b0EpPPDn1IpI+uI8kcXy48
H6egX1OxhcaLobBxrVjXKcBdvd5vHCLzYMdDLJASIEa65L1aiScP6rEDqgOcbh2OEr3UTisO51H2
/hxFuGkwU0626aocuYwIsV20vQ1MCUzKhFFTWPwGWaPNaIFWpsvW2GsaefFA1pDRrEY1ScmrE3sz
LNwO0GhSOXsNR63Ph44fxxnimJJTkuAMIkwnecSEi12NXjzsLwOv4EPqfawECOkxJP4qo2Xo2esG
rJ8MkPu2JTv2SY9FkDFi1D0H7QYTvF+aDY/LXKQsERkxzhFP4n6adcITp5h6MNEQT5jd8Yjp2DpB
KuRZaWkkcpt2mj7iNFmZDJKOv96CviK4Ps7ILhymCqsKAxeBXUUwl/0PdIPmsm6Aa8wSffj85IUS
nBF8ttJF1GHYk1Uici6ElsX5Uv6XX/kck8RYM4OoPwfG2bvzPWwAK1CbNLNeXXPbseamllY1yD0A
C1ZOTiqcJsEfGqo9BIckM5Td2H1w1CI07QzL720fTvSh4enxJvVzb356HZOO0umiW87RHf+xJRFp
QCS4JduCDY1dgDaGAf1zOUEL1egThT025KbqyIbhGaGtX7SAD76o1KhlaQD3etQfub54bJDAZxb2
amZAlTgkQxn6Mq4rr6+qGZYVzsnLX7+L+ZxgpL1pLyPZDR/T6NKHHqGh+es2l5FUdKAs9ysPC0sl
d83TKhPJQl8YO42l7YAtwFazCa/r9+gqlMIgFj8tS1uJY8etXyEtIfek2FG4AcaiFIuF4Yv8htFZ
wIZe350lPVisKb6D9mPdNNpc1x+MEE7N/TZyt0bDUwpoNOje3ZVExJm8hcXXXf5OoSZnAUkmdkZ+
6KW6x+d2ngY3fvN1ilWH/XMPDkWn/JLmL+Xt8uM4Rz20aTKozyG4qb+yvtYEHLSIicffO8lpyUVA
2L7sicdN4yGWcK6ipCS9/0s3lloTFi96GJUmxMoBHa+UYwBTnBWzVd8IdulWmDaOMXkXd9t2ld6I
geYLTJogMfa9Enqga5VR5gYBXQLnpWczNjc50Q7z4zruuW+Nygt8irJisCKY+eLj3FBPuoHYecNS
yHp6ddP7vFtsjo+6ybiiZUajKbCTnu/RBShM4K+vnTVctXIrIZTfdGXc66B1tcwJLvBeFTaGwM8q
hQklK9uYuTuNYFzN3XuGKqYa7xZ+7KtNPVGrw7uXOT46/3mLXVacwHWRjD1YsWt6Wo6ohaMosR8L
fPDpubtTtGpelyCyZWwOeiPVjz9U+rIOt0c1Xt/w4KIZXt0KxhKLjqvSyka1/eRnJBAb8y2fxCK/
ZMdzcZ82ureyIS1+CuxXY/K4h3ZU8He5Y3EcVoFWmUavhe+xpwvXBB2Fk4nC5kLbNV/GzwPpuxZT
AgXXMz0E2MYWPguYYuv41ggGN/SSgWq245VAMEIAUdATCLlneXVXxZB8HBDGfBfeq3hLo4VlIoUq
bst+of7UV51wzs4YsvxgqyRNcqvbZUeYt0Q25iGsROv6nK12JnDRYDX4mZnYyiBm6Kdn89QgfDh9
sGRlNkERTx94fHpF4U9uTEEZRIf116uQRyG7VC9plsrnCGy6XSXu1I7no0a2Fd/HeFBwJN6p62Zd
UzLZwrzYTcqcD/s8XQmV7YRZYzKTDzda7WTm+viK/eOPg9QNw6bioBgpw+mPo7phE3VutRY0IuVr
xPhjidIMHi6p0gW4RI3oUPpXCPKqae1zXxjdpoiIxhB0XsNph4NYuwlPaWudwSacvN0Fzm1KQ5R8
uPJChnqEy3e516etQBwtrwr7C82ai894+Sc8KIrpN36D1GFYP10+M436dzT4knx0/hNalqVokTTJ
2EeTxgg2qH3DeZvZLlJCIzQXZEIOjceSP3ZrljCREFiz/tNyhASK/7jsuE08IHxsyuaXYJH14nzx
tFXh2dLUihQA7OUpczuzZaTmqrap8zvNH0gYMTQjamYeXzKBeKOsqAKvPLhsRBNvSUy8eCs3YYpq
KyAdVEsuap/f74aL8oNlXuYP/kjJg4e4XXXe4mF0umlHwXIqBwg65iEsc9sY4qK00AfVnu4LzCVR
CjUr0E6Cqc4nm60//4KWbj9tLsvo1ySlQAruRtOXk8gpWqOihpW/iI3p1KS8V8jrfPGUsnZlDDrz
Ediq3CRWKrzgZErgpErvGabaU6IUg++llt4n51WhjJDS7IBqvGJlGy7+FqE8xu9LpzrGixatMiQ3
QsPr26etxgmzyN8yKNXPYbKDfOCacM5tNO+HxYjXfGq4oFC83oYhySHfwJXyp1TmMFWxGWAWGw6V
zvpgTTKhr2kqYJPn8JyhVHpwdL6GwfAsnm3+tobU1X4aXWI0sYqMs2PYVs0CjsRIfvx5JbmaoDMl
saGz7fvsQtzWrxsaChuFkSMqyDPsb9uX6Ew33hS9clF1KiwoPbfkocUpGMbaXu3RyIF884Kw9P4k
SQnBGYCj7yebTEBsAl6SVSt5H95mzgdHYH8o1e7CDlT2uPa2vXeghkiGukyZ9Wwk1JNw2XTnUGKL
4AOn1HzKGgZT6IKgahjL1TEVMmjq2TTCo9n6DLc+7zV4bh3/kCGN/Cl28CKbvuyw5oG8qsIimAkx
4bVySmLvt5JvKHOTe9jgHMebDs1ioIBD5HB1uvEqStAZTl50SlIWvtcGIyHczxsEtZ9fDBBgA+mb
w9pOvdtmC+gsDf4T51WWn0akHofXpQiC7q30PM/r7meDoTyGsQ6iWv68fsHD+vir/moNWqiIrhs7
+tC9XF+GX8k8EQYgDMs6IKR6DtG+8AIUY7aMIQs62h7ZbHoZd83qfgXoSm3T8XYkTmgl1Mh+GWCk
WQ9smgZ68BRsL2yIj66Y174vRaco6wEGUzSiYd0c0v+slmC59KjX6hVcjwcxCHz03tkNw0Miui3a
L9PmKTgxkRuTDZZ/gLoj5gVtGsOtpBrd/J0zrPsxrfCxVlnJ64vivitSM3nUK3moh/5gQ87JY1uH
ZpXDmWDie97QstuBsQuET+drV6j+Dudbf3F+JOc1itkIPWc7Qv86i6TpV3kyzngubOXQi97TTuj6
sHqISpGajPFdR3nol+U/tWUpQDwysiJEoeMARnCfEap7tou6E6UWXY5Xq2k+2VjnIfoUgGjL2ZF4
6nZGNXw40XW4unCYpuiOoO4PZLmU47vPUR5YnHNdiWDahSrbifTGOweNHTObfd6wfR+cO764ZwmL
nNbM4XucmLuZDvnugfjgEFVPOfNBmO41aMv9L21UyMlHk9lOPkGzp+7yMzGL3HFhl9a/UDP3G4Hf
HagEfg+H2GHX456f5XNisYecl8ydqF+DdXk535fXL+0N+E+uTv4Weozj/Y9iMSqEoZwX1J8F746i
hdCxbxxUT8fmqEc5G1gngJLjHEcYtKkLIa2Af9isYfzp3f4B1jPPK8MNnoQ/q6KefyXCqHVSK9KH
rqiowcuYnFc4pivaFGbTmpkp/L2Px9iGCK2pAIatt8Vfd0s/Q7L52Z1raW/GlpL2orWRFh6Y1BeQ
jxPw9heXuwi6ElYq88CIsPCjcnC4zIMacpOWSpvoK0UJLnfebGA8TrGiaoL0RRw9noEFoLGJMii1
QL2MqF7VnroEMng0h8EhzaEk85oSCMF+klLaIOXsUmMs0nCT5s+2uUSIR6Z5FjzmsMnQHjxW658N
yHEpanrO4alIJByfC8cvOoqldR94gcSq70YeBSB22dE1voPkGZxTWj5swo5WQLRhHRpYwEAdlAOa
7MuVshyAUquegtcQH/V3tItUkBW1kdgB9/GVTcT7rzAfUo7pOcd0/pB9zldzSuBI16O1w7JlRo19
zxJsEgLbf0gKQNflpH8oEsnyRyPBbrdICGUPYRtNYztMrAjhSqebsCG+2WOZqBPWcsxMF0Os4uhD
MM/DmzDrSQRQdeihkKTMS38TiZjRjeOrTHeyd+88iQf5dbBPb7GVQ5jTqeF8ZEY6mc77sMSE44Fj
kk4B9m8YfijLBQCeikpbCjvmzSF0ChLKSy9Qpb3ozCfpCSiB3eeGwFe+rL7YOlv7KxtRTzuIGQhn
iDCJISdixePs3Og3tzz/LHjrCFCKAmsPWiivSxItpI8wFTjL6cfZvmJbGOrdBnI0Zg/3JgtljdVl
xOex8x86sytNedsh9oQYpl36eRRJul2SRoNw7TNPd8SttewGnzUQst5xCXiJN68U4RvkThMNwqMo
MD57fC9sAfTilZ8JZIvlSJl+1vx53rzHRmRvJbWnWRkIHr1SVU6mrRwawenzO8ix6X+9gu/znpbo
w0lF6mbqYJseI6mxWcMczTgl4y0h34PKJmykrzPnzpwpB/U0iZqvbS1eY9KXstRxTRiP0SIeXJHa
cuIjRtToZSanViHu6wmqIPlPwpucBMWMVugAKft24vhAY9bss3WygS9F8f6ye4x2afDcQhdnkfoo
+KjOe/3DnuxYkmOnAIcRcjfu1Dsz8rwdqPlt4TKczTYLhfyl4j8yfSYYnxEHb/UyxYIRKrG2tH4h
NnlLX0lK+qecVEgi8DasMCgzSHfK8DoZrwzLNdgisTBWuTiG50WS4dZtygGHyKDs12FsKIr1GVYi
Z+1/epZA0lr1VHU4gqQMBklvZr1KvrKC2+3CRTRf9xKxEST+uaDDPl6qVB7v6yu0C3/z38EqDaC0
6n97sjDtXLkSJkyeTCAmALKIm1HLrTSziHwiuINPdxw1rXlwQ2HwjPUmua2kwvZePPQbatsRLtig
BCIfj/W4cKv4ifsaZIhbhjc7tobi24Z4n9GIp6qOzBIsYUIUZPkyC4Q9/yCQ2u39nnSXLd78EpaI
3YzE7vgKp6mTL5xxaDC81utR94Eeov1aCgxFHVuxcuv8giZTmdqe5p7FReQOZqRTml+nQYHEVamp
ew7N0gl2FLRX8rWVD15ASvN3HvVT374y6piRl7y/WG7uGoubnoa69jcEMHWWUvYdJACzxZ0OUggn
TaKje9XquCKEk//paRNbTXaF+7dyWFrHBhwcV92Zl4xVUuDzTHq7QCurpQZFoJV/onGgiHZNGJ1P
bVq3Oxrkgp5FgYGzjFVNldzNn8xtPpi7DzaquaSlcsx5JFxhzdcPlsp65Sgfws+/wW9KWqxNclk8
OEos0ghiT2ucMfHWh7k6Vixq/Ffd7FEUYnEfd4bq0fIOgC+O/lJ0c+RlhjtjlWshfKKNt/Iga3Er
aFYcEQU1F7uMNSBRkKJx6pU68D2naFw5emVwCg0P9svnkssKuOLqsmEsGWLNCE+9CpwUmTAYMQ6N
AQazePql0XH6KKRe2UzcRfqvWfJCqHE60qEfkiZiMVGVg4kGta0JMWnbcAUd8ZWDh7ZhKAvjfAQm
HvrZA0UBJRUovYEMUG1OdHQhPYYXl6fvZ6BklsJeLUb1yZdVYtbp4JPB8xJ9lOaLZbba+vsia2dN
zEq6yNTWLN8BM5Oyh3Tr71/aVn05amLOhoCYDqpymZjDb+yeSDXB60WscWif4UxNmb0ltgVSWI8p
kR/RPAZqXDS8PYvbKmRdD1Xgemk9hNgkEVfTi3R8QRvScZNL1Pr6/AbbMVSyE7d0iCwB9I2/2CPU
PAEC0ojEdzSppqY+lXR5KzUhNpQIuKuRdasn1hX6Qufj552L2tEVfSOpRNw1AvvG9k3x1edJPweF
Fup7jggi219cEsCFoN1gMFGtV3BkI+9lHmPSOvg4QoIrKqFjK4q8ZArLW2bfk3+AR/FIqNSgBb21
XSmITGRUHxeQtcYWWHwRxeeJrCFSuN0qkHZqmRo1R138Lb7+XL9Y1QrV8ARaWh3W0ZR5JQeaWTsZ
WfJ9Sq4ZKBd/Tq1K5GYZxRPeYUdi78Oq5x9hQcoH7boPdsUxj9ibs3AUM/SB+EJRJPZS620OTFBi
knDilBibOqELj16rWsJDM4w/z6Ds7BRDeKJpWprIXQXKeU+B8PCGQONKVPLyfPsKs056D2VyzLw+
TYA6BPzr3akpEizzotWlAv3oVVfAqTZJA/Du7WDz6/nBon8aeZqdYazZ7dH8dDNvhx/GW7D5cekT
m5HrmZ1/96o2tWQWlibj7sS/E64TEotskFH1uJfFAdDXVoJI2sZQac4dtoCOEO3ZWDdXfJnWqvjc
8SATZJk/c+3h3ThLz/23On6H7fG+fzPZliRznqGJ1DvV2p5xKwmTaysKZ0r6+2+DS3tYZUhY/j5D
Li5Zy8kvJXUTZaJAvy1QMzg9yHnQ7z8gwj6NGW9U2L/IDfi0Yvq0Kr8W0A7q7pBHeFpTSe33IlhL
jmvvufHJiDMQtU+pelGX3E33ConkbzoixqBHR2e6F5ZoFrsLlGQjgsdDfmDLJJ0MlI1V9cXLcyzb
U8pjWh32Kwpzn8LEr0uEkq8dvJRTBsnV1mOD4FOWTLe0KZfYBJEatZOUkl6W7bqUCAjY9nnJG2cg
KygMbnzCX4rWiwYvXF2yr1aIjf5dlEkrF+7mvZRZosNwkNLqLn43ZFRyrSdgigb5K37qdQ7U2lFa
UbM4IVOSNusd58g8Ovf6bWfl2tbl4RlUiuA7WJ0BHLrJta0ElRju22wxfwjHmm20vuZBQUnq7Awn
izn15F/qfChKjkGzPPo9rFNf5J7W4tLC8HN1u0J2GFDXBWh12qBmIYavqH5TjLgcC/V6Q/Qlr6F4
FiQenijrKEJ9rr4/jKsHrJ5IsfGA2SGiFWBeszecrtzdwOZqCuG2Q2mOVkeetRdhxfDVGY4DG1U6
p76NsSz666vByoSFlgYUgzEeWo614m49e0jCxGsR2WokiWH/S9a7fAHuCo8xB0Hus25yvIQavlAp
2DQpxRXAjAVbEsDq+O4pTmccigiBuQjxYD1lgcC36WepSgrohVC1990+7upntPLnSnRGEs4spYwi
gFpUelKseOdQsSDjxzKBN8aEI8MjGgDFpLK/U8nPpk0J85tVMCY+Ktc18HPcVGwDITlrZpWYPVFF
pBnuttbsD4mKeKc3cahuIx5GgU31jNxHj44P1RaNPNjliipTkOtV3ATJ4rua/bhvPiiu1E2ok2ra
9kC9XDos2i/AnqCzDkGK9ssKYLbNeaRjRpbEGEq1NROrCh4vsD2a/rmzCoPBgcpT54kLMyM5FpF9
z7EC+iaYKYFQ3zl4FawCwgxwp9rH/3Fh+7fTgqcHje3bgd3SbGUT/9OdvReo6px/skvpPDp9NTDC
GbFhH5VrwY6ad5bQw0BBv+8DFl/0Mxd+xmpo6gUfoKDTDKxUnCw10pSWUTY/JyywDvFs6p99h367
T6C/OUaCPe/GaBMuW/CyVz+vUDMv9SzwCl8MFRPy+LTJvk06Y3LpETKHngVzZkyO+ueP01HlJum1
oR6/wGma7dG1ofMNSUpNcZA5D59iKxYPDy7ZhJfVoIu3sJKFMsY4LgkohBDfthPFC5NxpL0QivGS
Ct29CybU+3MPR56dUwRuX/tu+IvUcFlMdxI6Z5c+jFUJwCW99XBoiHqFhAIlck7ARBMuCxJgCKV4
mKYi/GkuFy53YRjC1nJmWbHR37jHea+9MLbkFTcs9+wt7TGLxO/wC5xwxaPX9Ta6AYCOfHonSTh/
kJJFoj7ym9JurM4y2M19CCp9PyQbwVCXZsq0JNoFh9XKJMOZMr/nuY97+nNlPXZY5cWCzjKPtpN2
QOIdglTJgyLC+pgedoxo+Uqc+XTQiZh/ygtCfY4+Sxi9b5LIvBkgmggOiTUyBOk1tfCjIqDaAMZD
lkaEbJ8Kh4qx/7YbQdddTVh3SpLaqeYrbgnF0OgUETddr6gbprXvdq8qO56dCRORaj/XTIoq8K2Z
sfWaapE5pNIdw/0R/WEvHTHwFJ2XGzlXosIH+5X9tFbF764RSpEOFHgaoi93l6n+eUo4O64OvttE
tJvgSFb1lv4ztXcVEVAm8tvj/M+IbRDLy2FYXkm1tTjGH+dcuxw/5Ov7/+1L2g6iSa74THJCR0Mu
wABRgOPDn3tkRvz1Kv+go2sXjtaNYsLvBF1glx4Zx5TaLeIAA7L8j2apa2vEb3lReJSGQR81fDKl
7qKy7Zy9P9hJMFWU9j7UXCtonyYQWQMfCa01cwGCj1sZ7eU8jiEWxI468p5xjWH2gwlDiOmDIqt9
ZZdgTqSaetmesJsU8IlOXYOgHrkkTgyX1wr7oWqTxZzQSEyq8Iv4C/HBuqF6f55KNU8jfprzyPWI
iRwUNZSWKhGtT3sLA3FArIExFCHuEVNjMhD5uDr0muP88mltwcflEtdL+PdUNFbBgN6xf0nxzwcF
SYNXKHpsiZ0+Ihn4USsTLxrwdgUWrjnoN94FOWaa5TxPMoEIGJHbsbPH7xGfhwcEhaPNlkXIyldC
ShENldku7v/zb7srxhBjD94cYqlXrofBHXi/DZHVcFWA77mRYLEZstuGgDlnNrqc4NneAdUC7XK4
IkIYCV2wuF5KVC2ksPof2QHX/dgaGUF6TELXKc9Fgr4yQ440bFUWYbNNaKQJ7ak+UxzUteze3Mh6
LmtVrTFjG3G3NKuMCUrhV29GRW+s4dF+Yxu85prVakydZ8JrCXK8HIOOI66oPg4vc7HM9yB947rr
Tzirrpk9F23zjPrWY7DrnnXV2+KV48xj0fPDdtyqjIt5mSxkVaCgGNPY0rIa670zmnAD/54ZGJ4n
fl7W5jYvtqQ4Uq6lny9bYKmBYjSOolmEgS/gc6AyHMHG4pjbry5rdo6vnbLC6THdT8yhY8k4iqua
4OtUQPNSJvF/tBp6ewR2+g+pHmW0Vcmphdx+Xyg0DN6QzNKxs7KU5g++D44D7iWzhOilt8nI7rP5
f2ZKUW2ERVvrkVeQe2VA/FpGPrT/l+kRL6hfU87Q1hF6i0hsu094+jtAb/pXCKODqde+UQ8kNbcA
VANHR08oaZelhS7gTEdghEfg2XecgDvp9TcTIrQz7gFMahdOw3UyWsQoHK6mKNhUR/cLvMhdkFJi
vv5l2XK+I1CcUrG4O/Qi5mARDzDDqzV7YeoYNPpNSHOTcCqJDXWtcnzODxmGem1Fw/WUfT/5K2zo
v8lJYWJt/347x0i4IIuefVsuuAuXumHQbXoabO+B9MRboJvbkK++juAESoVIejpPhKw6sFsVl5UG
5KULIMO01/beBkY4T8IIkf5FzluiLqPQI/EeNY3Sq7tIrojeXBf19b1pyNCiMGfovGSbniepijFe
YsK9GgphXUbcrc8xEqHS3SDMX5idSeCkDkzufY18zuGMeqkOcLLu2C8LArn3LoGQxyKCV96NGXyb
7XkT4TZPv0+M5qzt+QneKkNqiOHbQvfjlLNwK9YdPUiNYoDEPYSIqbTS+hN2rg+jzepIxeUFbfSB
7NGxYlkoZSymEWICvyr1qi5flJpzlXGMEJLHTNfZZHY7py8zBnIJ/9ypzP3Gn4KD7C1NmLO9mKgH
bmH2QzyyQLQVaWZ7dtWGvf9Lv8zdMsiIkcDJIQagGorQ5cszKGdhyNURq18uf0Rg1Nk5resQaCBH
Di3uk6/y/ypICqBWQ7ghY50XfcrDPMfr1YQKMp2Hj3mUNCYV8L25LksiGwP/oL/T0/k6ZLBHec7e
HPFY76d1R9/YlXWIOIWJejGqabdZMHqHniLdVLT1T4buFp1ShxVk1Y7kWSAYoVD84CKH9pd1El3Y
FMvVV0neDUnNaDBCtaZ8nf1Njstr+qF55O25fUvJtgThOmjYG+qWb7EVt5sTCQEUnRIJ9dpQxG2g
l9IEc4kdsdoESLOUQE9mYCoJyniJgAgL8DCFMsql9n7LeAt0Oi4/UzgObCoqVxqBk6haRNToBwxw
hwSPAcGs29VjWSExq/V3md0+HskaW0qgC9/SydYib6VnpmMSNhRuUB7tGuVLY2qyVRzZcCRKE4Jy
785JpKRm0u2aTLWKvFFX6mR3igdXottQoNIklKvQg5NOtQ5tk3w8RezgSspF6cnmwCxVj/6HA7gO
k9kY3A7xZKdSulePrl0eyw7U37wWU4DqhktvZN3cSdGxj1r0mr3tFGFl4rtY1E6kpOPJNCJF40v7
r5wOmD2Y4gUxk+vds7eu2S6gO+hRr1vhbEwueuLJ118lLi3ntxRexg2CdqZZW6dZk2o/W5BEZKKV
6uUcp3+GSZyYl4Sv3c9Z02W3H6aGjSs0jDWpXdSk2aCzTejnowcEwHkV7wh6owAOHOrTebPWIOAs
Au7leXXIoiIg5uNNt1FV6zkCF9wAPXAkB4fZQVCFTUgfCGQu0XO1XAT80eRdswUdn/zIez/2RMe+
yeIUQ+dCzKqO4v0t63vX2W5mMQ8igyccMHHNEsKL4NdlJ1kPJ25Np/5kdVZsRVnU4XyxjQl0J3s6
7ro117t1RmrccCzCpLbZrQV5wl8jF1PLHrxBoR6lLiNXeGPveoxt24K2z7NOeEZcfMemFQtUbS/u
yW7sW8spb4sD5bG8cKeR+AkpKP4pI+ZnDlSM+JYcW8Mea5OrTtk4NsoGTIyV6zHnbWtW0uupM40E
cIW0ZGteXfnUwPh6dO3c8gGc6vJUeLxkaZ7ObUfBKj7D0SGJtaJlBykNmLd/8Ux1HkGZNMqO/wu5
4KhfO5ao4oEaC2nOuIiYi7Wq6Aye0sOs0DGNioDm/CFdCU181AwCyp/oEp4gTdQPtzkE0lmDhYhZ
cey7aOJ9QgtMsnk/UC4tI5xDU/rLqyEzZXAjnvyWMoaRelS+jJEPMaLRXNMeDeXuAABF/BrZjazS
TV8ZQBWYwr+4GX8owliPr2uNJQCMLKz0eUDD7iy7x9ADcr0fVpqCPALX1PsiGwam4F3yfKiAOSqk
chuz+W3pqMHSS6j2GhxSaqiEqESgUoAbLi3fXHhLElqYRT+NPU1lkY+Sb2oUhpgcsRyPPoosmuNL
g0lE38+6v6pqlmqxOHxFJjwtTwDJHvweYU+pGHQ17hDiZ+K/QvjEPg0njYQ3ZOidlTUyickNscYl
Muyo2AEPQ67EwEaiRd2+HQm4ud43nEMYUVs5XbqqYenxl1AtmEej3nTzt6FxbvhI6N6R2dcsHnHD
INd7yRPHpUap4icDrE7IkNuuFe4qwewsOatd6m3nuzFMSWraezvgnwfodJoYCPfDblVAJ8CHxS06
WpTux1xBbNOV5OYc5DZtTvUI8K2n1X3NyQnUqIeEsM9Hw8oNec4ATxeFXqPt7zlGpYInhSnpyQy6
fRBz2KrtGhSISm6/i6dEOu6jrO2aWvkhFK01EFcMYI+13SJnMaTsCQvGu1vbT5KKCyoPuUDq3J94
+0qI8huZmEzPTsj9Xs3pPMgLyDStmpPsRWPbwV3STtPNavgZop+rFg+z4/cQm2vkWl+XC9aYX4Bu
K55ZiLQufgWrHj6hIBwmEVIhZwG5xl6Zi5dJr9a4B7+p6StiQS7j0v9YVMqrlURzMWgIehGwq3GU
V6uNTjnZk3Uq2fes2aJOcxehXn3EskKI6I9P7+pohwO53DCT71RCmG6GYgCKOU8jEmYMrSlnk3ej
IZ2g6GgG1D3mX53PUOWEf+f6OUg9thoR06yml+G9W/gM+cphWOt5xXDfL2FJnnaN7dBRm06Tn4Kk
z1GEbR0ah/Y0vkBgZxt9YAOL23i/4X8Egy8MOINMaFqADTv6nhwA4YPCDGnezXsjAkUDSF9zlDmB
e4u64UKDjC2QQvSxpn2p6mq0U/gThdH0YuJWr8522RiiInd7CeHYD1/qZV3zn5xRP4oebqA5WrQW
bBBcRIeyz7eYqDnw4awu/HwdJbiVHAO281wwRjSi2XpICPMC1zxndObjYudPRA+7tPQBwzZH5YCe
CiwHTiCZowW1zcni8E0kGtJGo5XrSNIj7HEcO9q+iddFUxRRGS4nvEnKMp8sbHn4QqYJaKntXD2p
Do9en6d/eY67xJsSMjxkj2yx7EqyJLzmYT/zqiTT1EV5b1lypRrZYdkpFc1gKb7l3RoQw/xZsa5r
DIE/5Roc9iFr22vvp+/+Q1CENsawCkirlAMYiGzK3Fy4ztqUHHgHRB5twKC1QStiSo62E6XVISUm
WnPVJxGJWNNOG0pw3hduP1fjbV1ZnwCsslvKEBcZ8w6LQjd4D5vTLVvr1wiGi6/r9CPVtEflXItt
IS2eFb8tqwBRwky6xb1NlooU6oyvw89sdqhicVxBW4SdpZcIsYVR0kSGknx/A9W1T8APuJo54T/1
0wMFAyA8UNwtAoFR7gLaH+a0Bsfg1gNVlSx9vA2/XDBx7QI12afCL9rmzC+qBh6XRijsMW7Aq1Yv
NuC06YsK1YKAjCJoVT0uRyKIbiy/IMYY9r+7mqTcdzwr375d6JThBymDT9dhyPpokBRV+OjDvuAK
THw0M/pjNrfXweNJY5yakM2lkV+0nuX1hKQ53UNY7/ppODm8xzIEy9mQOUF/dpyI6j2PskvraiUO
ApkA/BWp3umomJfyBja62ANcVcYEyKCLEriX/AFuBSGngKJsDKlGAiy9yfvXkjZTHH3q+nZtHboI
s8nX7MCVn9UgcLjG4jKP1GmO12urfSAIGRiFia/pQAC5St6f4h26gXIM0nkFonQ54fZpjEOZ8uAB
q7PdZUXcebxgONoBmD8ya8bCYGR9zKIksWHu70qNYhyQ8X5MAtDoTC0Lk96TXyByGujoppbyEfSr
1pfd2F+avx8/DvLhXNdVQG1lVnYu3Q4No5z61bidlf47dSOZnDieEI34xCGEZGm7207MP4pckw5D
CyywwaddPHe3siJeBoaMfEI71TBcqyMlIglcG29nd1TztTinphMeOjgkcdLyJIST/NVcEF/4VU9y
eMpSLov/9CxzgZVQ8YOiuBlOb+irCuzCYsHm1l1MUE9QlhCgxi2EM7KOqC1qip/Fsg7CZHtCkO7G
OAxTJskjq+1rfY1rVGug3Gh0g4idKMcJ7JfXBxmXcdrCdzt+OTQD+4pG3Z8ICmb4dp9Kd6alN3Pk
GUXEHYXikR/sZdGUx0gDgU4ocQIgDm5WvhdeRqs8oXHMveuOfSMnpP0hTKd56qHvRqWMJD0l4dvg
f4MtVMhWkg0uJklnbncWmAG89oWjjsOE8iEelUe/fmn3YvM1ZtUM7CGPUyC11SighRjWOzEn+1OD
2x5jdj9982v9qmkUInF9jHeMMG3xCe5qoLiu0hUYR5/1b/B2w4m94PbrfRc5iQTMG9JRXgdy+J00
iEWIkYGSreO+k0BUf9FEphRWeJZXzvqzxvY7pxfSuCLuyjdX2BdIFKFECuKEYy9WJKD+LZRnl4/W
qhbvmDiO3vrwyoVkRDFz2x5WfWbEzqJ9LdDMwotWtQGICpFVsyO94yYT3h5J8Z8CVhU35K7L0Aeh
/W9laRPeAsDb+oi8aYw8mEgCuEwsw2roPZ4XfHy1erLhQef7nsj3noTXTZShRO7OhKjgZF0Ocsvf
J9tMa7g4vGGz8SlDZoZ+EWA/Ss3/G6XCfQRXMlOiFvs731xl6rIMnaQeU4Q9ES+duzEmR6YeFcvy
Nm0J64eMK3JBba+9OvzqWO2z0Ne9GzyM2AchHlZcDmi8ShO8SkkeQuxuOTJy6OKYZEGnSSGS/yPp
w2IfISpnq9L/OwO4GJhcGVFuRDxinA1065x199wmZgI+uG0yhWQggVpa0ZtOHUiczIoNgJ5znW6t
nKCATRjKwvAEjciOjyd3Xv5ym0omkB2znSCCV4ts3kLaTwNuF8wfLOFrXWRp06ZRPQqZ0RpdvHtN
bccR/fMEAvfisCETUnax+w6r3Tx9nCXSIKWkADVV9EUOQKbbHpGWjHnnVHg45lNEDf4jcMqL2eyN
DdkDgPbkU3Tf5bSSwVZh7zo3K8qulL54tpOExv0cgndnb48ClsKaMcHQGfkCbDutD+BonVvtTTzJ
Hh8r9Pu6NfqhhBDy0GgJksSY968m+wvoQM3tFww10x8L5LTcEwKyyPpVfn1KDCUCwIbsxLhyTgHp
D8EkdKuX5okSa0FljahabFJCbz2TCsB/YATaWP4xH85Fe3NoAIJ1jW1OrbRpwFyox4T2/a6DlDxn
fxXkSqsuXK/fwShxHLPPMCuARaLd0D8J+pobX3IFo9rlL6OTJzKdzRmW4xXiNx8jTBgpWWDbK9+I
fR50Hhc+LPzlKN5iG4F/NbK2R0f8PWjlnu7BJHvwiklix7jfg5wtVn2rfjnuAjjb2hfiFoahzftE
EQMW7tddlqAfpVnj8gt1VYqky4v4mxyMVVyUYMVgwc0MKSjPmZ0GwN9sZcZVH+6J2H86/+Hx0v4f
S/oiDdUMhOpdksGH6zq0vF5HbVB1psVK8/GMAwszZryWsPrDkHsKExKzGGkBlclAI4EUFXJsBspQ
ElzJsvjYKSoUxFL9fZ+h3VSA8fOoPsVpg4T2nKLp36T62qjk8HpuYYhEEMz3UfFoG3vFzc1/CeBB
ukH8neHCjw9IsAMj+SpAIsuA90OoT3CgI2wGWEpWyY8Szy2TPAM8mf02qkC/SZ6RRfsym7H9sMMi
voJFYRzBqQX4kLvcMEMMU0CrK/O6LA73UoEUQRi2Gqu8Om7DYogMsGRsIzfbGwOLZ2S7LYvJriE7
Eytzmlw5fJB5uD+e3pFgGEwXgUQ2GlC2smj3imc+dH7Fht0m6UNq+/DjqBd5GmhRpputUqUZI7Ig
rp8MIEXCHHfP9bvZ+PGHgAM+WTMlt5vk/9YZDST6BGvPRajnBnsh0Us3+lHu4cd7laU0ko9T43tP
MZ8SpxEfQjiUSZUd62iaIP3vZHiBSRacs4PGHpY9dPJVqi320wxo5EbYS05u7hX5UOnlZ8CEZ7oO
mYjrlhfD8k/PAKpeMf02bJWGP3OyUwTVjVqzM663agrm7Ee0sEVgBrBLix8PEqXyNYe0Q0EaQmRs
A2ij61nhsItumVKs6NT8AZzKPIHT7Rtfqy/io6KMBwaZQ9fUUHOyTfIqib3e6gGvhkKXezDmfrir
A3A72czM1/jQFeeTTkHqnceW8rS1McdPV+X2Il3IDbdszZVWGd1/jx4UV6ECQKoSwNI2/C1Ncqq1
5ZZXzQtbZ+ykLdEtSVzkMmwxrh2+WV/qo77QJzoCJRo7hw3V/otRywcjQX5avqCRZF4VmuvOj56/
iW7+4XzAG4tm6sf9borVZjg28t3KuBiT+3emsqc4m4vTBzS9rgHxPyALFYrGggmFjReG57W29BNs
BgYICwIZoDIr+6w/qJ/iErwRHf4Q3F+7gX/DFQJbPifKfm3kwZOpXUfrpDiutA390TcT/II8VM93
RAlhN7oxh9HXL5sIg9tQgOrVd6Cv02ev9/p/652RJ6S4MifJN9thlO2Z155Sw58yz/CFGKM22W56
1bgGt+WgXoFkpzkFP4vzUYjTkRCkCJcrJwSsfN4ixrd98OBS9WJr3KYt7YlxOk0k24didFXdaVuU
osIrqio7LKGFF2nub18AWIeVrMWug8w0ook6sikQ1vXq/CQp8nzF8ARX8iGX0R7U1ketXWr+rHIk
k+mrrxz4Pwxobcm6eIwGArfR6GVqIRxM49QBreME2bexXoSCyW6KSwtbHavZ8ocmgbbMShfEPB4s
emgVbzjlvHIo+oB7m9R6VGYbf0Qz2rMDozKAsrzXUQgBf0Qxjo6Nne3niykDjECw6NlDsoFdaBOL
4YEzYOo8MdvAUxXcZvJc73BNSinGW5WK6qX1t2b+yWqALTZ7y6zGRsORYJpsQoNF4YSs0KzYimyH
Kzn6Zmj/CzbXV/MigH8QQZHWgsknAw+6fD4VFFfIerDE3i/I7dWnj7ib2DyGVygdjAEJ1TaydxAN
RqhAWP5Ie2GllmGJnaGvNwiHLascLYXYaAHY1yMfwaUC6GkmBXybPElGsmbPFOcSq3nw1WnTxsju
QjhyIREIaCl/62uEFE1aixD46HwVqCwY9z7dtrFvRXS4rPIGLLjMkhQhVCdEcBXLTf/McJju2hPh
wUZvfM2KfhBETCXJmqx1UIT/bZohBQOE4ll8KXPsFOUnC0qsm0779lYRuqyiWyQOqZ9uXPM7DcVh
NMmci3pQfW+VDYrtwNsGZ3xe7Fb5LGzpMhIKZTfCG/bJ7I87G1feU9ocHUQsWqpGMgvyy/Xx7i+t
+NY3JNseqbboGyRXCjqsnyZ9VK2hxbP3M2Kpv/jP8aMjk5d21oLTWXzkWUzGpDoHE+Ss9b2stgaE
aVuu5gErj9SLuU2zq73B2A2mTH5+p/vySracRnCy2uPsO/rNpdkcjxH0pUj9NHjkV1PoxwYWWb8o
m0CFjUbvx0dXxAoPDAsCwM2UPl7laWaICYBglz9JNU/hB6plIzjyOI/NMBk7eQ1h5RvhA0VxdJr6
wuca6k11wORDQ6CSbO/d5FYB26gBCCeMqd+LWUaEs/jrIH/lOboOz924xImFlS3cS2Q4OnsahSng
w3+dLqLGc7/b5XU9A2sJHby4F/XQxGEkGWqv20ZUCqsm+uVHsVR96Gm0upMiLOOnXg38P7Adm9oj
gXjvaZqPGRELfbnG7OCfDziiears7GR+za5gqIgs+Hrm1IvSIjX0EmWtXwpfiX0kygPzWrpfN7Nn
SJO4a3jc0v3cjPeksVuu+vVp5BzifGT5TgLxX7LloP/p4wiLQiGMMa0cDaQ0uW4Nd2n7hdWiVpcr
ziKkx5qAUxpVwjybpr/8Saj6oQOeuUbkQbMce1vaWtxFj9w6Os9Is80YP/h1oNNgstvkGkQ7BWnL
8i9eyo/GzEpVnnYmxz32i10YwpkMj+tYmE+cUj/xXGXxXeBBKvGkN+Zko1hwZiaat0l9gwkdxaTl
1VNszaxoLEM7txNfb1PO2XyxEtgxrvVl6Hk7m5y1v7TpYskctJXPAJthSubXqS8vlQMk41rXy9UT
sQh7SKQo9j1vVfR7+LXWsdT0WJYJP/sKHBtrU+1hvtvUb8Qo7RRIlpaaEGqaqqARh0BfUsL45RB8
d7/aiORgTcQepS5Ge3aGK7dfPfTRPAaPrh8WT5YsL8pb5uyMa7QnfK8laOCzb0mBUzvwpYUWjk7O
wi1dezb3lySdRb8a4J6IVtOHaJmw+diOA/1b1VPIEiA1+Q1UyvPDLpEEFPFFImVTkKlJqIgWvgl6
NPnvvfzhLC9+1IhitDqQ7J3qTAfdqu3XdWuEvfufIAPX4L6Yegyoa8MGKIqABnJnjW+h2HQJhhUm
NpaQyLM/u7qUGgpzFiiKN1RwWb6WW+Vv1+aYJvCVN29d3W0r/9OOv3Vt+q18ETQpHY0Liz13yYNr
ZYy7jeFegUtHsbfTLSTcSHqiFR5ko2weXaASAFjaJiJBT5bPBkblpExRZuW609ZokRAqmRrRCJK1
0erUOLNMS0oBB1iY/oRuC39VkdWnIZ/J+C9KC6glwPWiEOSy2ACxFtA+AZMKKttMPK5JvW9Htq7I
676/8Mewoa9KlWXFg+5BHjftnvzRNJEGaxVIyYof6LX2N6fky+nbegTL9ijml/nIeVv9virumHhy
tC1sI/Tx3SK8wA8SK/HDywmwnwZk0I9yiqEIcmDeQLUA4wE+bM3ZNWJBa+XibcDE+Ltigc+qCYfJ
lC+n8CyPX9HdM8GueHxQi8X9DMdDrsFzc4+bi0A7WSRqEOR/xIw8B1KWmBw0x9jMXFE8BX7YQHq3
qOhAi9cIhv51VImmlyGaLy6rfQ2jXa26pgRhF+pJv/zQxilgQJrCyc8YiMeZ0nOmC26SQTnRnnKV
FgS59ianCyFoedJ0HmDyN9jFjTu3v5EO0FwBvCbg7oHgkkEyYsOvkSYTomKEoxlNkB5e4YkxIJy1
41TO0Jv83geo/KhC4dc/BueA6kEpQOhA2r40WkFjDI3fOmPtrY4RrsZ+WHsp1DeUmkOrsXw8UyKI
0l+v6xfWlo9WA2AJePyy5fZ5meRQM/VVsy2ymYFOSNhIJVMEq5mwLB5RqE24f5/bqmINaE8qXL3h
rIOMuGUs/CKMW+baMwpJrVEbXe5yxH3Wfs3QwBDYl/Yiqn0bDA8J2yPNLwlEWlemONiHM8Oa3tk+
ETPFklo7ESq4eIVwSEmVfIDUIqp8cWCfrXg2vZTYVrcdrXcwOKakRPe096Hjr59KH8i8vo9skySx
770P0+b85BLsO57w9HBX7Mnu49PiT7zMmjjvG5ngq9JAdhe/euSkshI/X/q0EbPRDpESfO8FU3CC
kGCZxA10dhIVoENP5UPibSH8+UDoHOivmOYPS6mZG7Q5hqC/ILkIKIn5JVHB4IkRVhvsVqZP7pR5
+IwwSA3n2JJ9UjiMvR+ZTl/ehfLZyrbY5H0dzP5caH124mGYZgawrz27TxbewzXBUcfDHGM+HVpi
1/fizxiE77QGmnPKNe4/aIuRk8CBIeP9OK5h4AoqUWSwybUJIwPtgGVp7iThK7tevQ3n0gy94Td8
HgxD6HLT7ZflgIun5STSU8qiA0xLNusWUrawkftlahBvB+c9D60rLKXzjYMwR02LK/wGhSJfg/Rt
EjxQpGdjBxiCanPqqzTzN20BfqvqwW6fetMYEff+1cu3xCuVwjOz56mSVPuVhEx3PC27OU/Adpg5
C0bd7svpa7JOPGCO1tzD9xCzjK8aL26SMR3xC7fJr/ievuEJFWxesJeQ1eR86kZNtph/Wstc+UH/
pbXSvV+uKGyv0cm96/r8bFblP4b2/aYjQ1jpcu5jVpWQjfie0v/03IrV+xt5ecXZepsbTBV1atSX
pP9Y4Via5LrEgbCGVw8zrj4Xr5Yzypvxt+tMPrJivQgLdfiBCL10EM4+9oOVE6ixzttpvZ0gslRV
GwwTUvjT0Nm96CwkINse+lDKqd8/5GEx42RSI7zN8RCfhy+MI+nZw1+a927HWxYIg7BfwsCAUQIO
c7XNCtZ/qr74CrCLLIl/SXUu1FAx2lKfZBSCOaRwO00X0tECsB6ArxUzntl8kCVcbcQ1ktlHXl46
bCiaxZYY+6pILvqF1Do6/OE1gIpmztOCtT330bTXnt9Xeu5GvJP3nzeglE+CS/ve9dr6k8pkHljk
D+SCGsnh97lpTdD6luKXl/H8ti78wIQ08rzX/cor8ww9q8huepoPxme870o9g/HGTAwma7fviJlR
SmlnQ5+z8HtUyjDO+GI3cYQe7lS0nWlqAkbjjF0GxIbk8KX6bfQqfJ2v9Hg9BOG1YHQ2YBU1Vw+w
vYtmuSTsiFms4A6rj+tWoBLN8FqLcpj5bU1TYKIr74rTWV3yBWXE7JYIzzCn/4zUYUzfP+NXRUvK
Ukqz8YvUqr4bT4pKIsz6y5/OpulEBQxBvUNkr6se4D/bNjWRMVdW49vV5BF4WTGaHERgRyOVv0Y2
ziqfJM4ok8QQG593O45hS3fapjcxv+A/+CofXtmr6Ufst2S+mQByk3/ngX66V7lrbu643MIHLLxT
1hQJ2gbOrKiJwHIeQVjlEXHTzo3oBrUGx+WkGVKa/Hjqg70KPqTBVexXSBNrbxe7wSeCP8e//4cE
EGCCxCp5CIxFxC0zMcdUMcGsmZbq9TDNSodo/DnZ176rSjjBrPCGhZa8epoTFDpUi6d1jQi8WBmW
HuYSN89Focg2SBjJimnBSyy/go0ucOSaLq8wMyXgkLJPPfvDcGh0Mei65nEUjfnBB13y559F3IE2
j+UaH6h9ug6SDJP0t/sz8kgJ/cjaov/3CTninThuOLCNJXuUAvobeo7J5HP9/kWLftiFqjMkY7hf
BEI24UXqfsrzY5aZ3MPjYenVYIvZRAvbNtZGbg92nv+QRalXJv2vRkH+pi8LjyFaINeWdV6qRA+l
D5nYwG/+yTE0ymLCnpuGL8LyXTH9ik3QzOAltnlaWSAJMZrLyCtaJdOhTKR3kzLqZ3cJ8a+t95pl
bDSN8xcTwPIj8HE5nMTo03VYh7yOwIfWtNkc7vh6UgrGrYzdf/SWwYyZNlBjNY6JC36x6hMBNiXl
WsS1n9kPTTwPjb8qq1KpaFFI0/QuHfCSh8QIqfmYWizFRQkVYEXzuwHru87tiNLhle4QgPiStcoP
KVwSJEB19zjW2FwEMov2PeTyOKWFSTVg0jjOZgJ27CQ6IilBKwMHkWh3jJh+paSQQSB98RCsH7UX
572Wb0PuqBx0gjQBU3PI39i3L7LnM01qkvUPQfT3jY/T1YCSZb2lxR3tuPcpDnYhK6s1W74r1Rym
Zr5pmP8daAPIWnaFMGOAv7KM3Fi8gyAqihOfLPkywMvPhKPLO2lk8SlKFnRdTk9xvsSEYglIebc4
mb4gWven2Ktd994ktwoPdLx6pJfMoK4feuAalmL4v71y/OfpWVI9Tnukdk/QsxPZNsmvZA0HO32C
SXrS9A4irDyhkLBpbmh1ZHpTpGYAhkGhKvWWD1GbxkC+pgJlPF8Y7G2lgOP7cR07rjWfJ5Nj1FVn
7bv4lKIo11+m0XZEjaIPiQMOOuMYFuJZbjKnEerczVeMhuAcJvV03Oi7Dq1z9Wofl8KnME1h2t7i
STADb1SIr4ym0SGbBOIanuYzgG89NPCMPt/9CIZci1/RAImcx36bNiFxz5mKCB4Dr1++7DnF6zb5
OsmC6DsXEqqMISQ6es1CE7aUjokl7UDBPD9aEIrZQ9SoWj8OSKZ8OGtYURq0OhFFfwdQm06bP92v
s9aACnccS4H04+FWLhYTaxfYIX/SIG9qjR114TrApAaC2/tJzEi8XJ9KAsyZu6aE5cMDcarIp8/R
RYzRZAJpB7+hVXQR05by9Gy9yoYYO6DAwE0FFUZXZ9/OuZi6c4ORisBpJe8kdqWC1VDQNgn3Mlps
degpt88b7dd6KbHCh3aubJmrWHWQ5XgL1Pxd6TDbdM3mtKoLHjhbzvytOoWL5R1cOqRyZ0j8Ytkw
ihj5/fitJqQjRTbfHYoJGukeCdNYXCj3qOg5DVUngaZv3A6iojwCKONkHrUQMTxDLDsDuWKKkuLq
fD/kEwRFaLSimQ3dMa0bFFUWE72+XOVohr/660VknwrCbMmDZO7XHjrF/h69EpT6+U32J2pIyrPL
jGYCgnib2VxMFbVr0+f5j0DJ2mI0vzcF1Z3zevwjmJfCpRm0mabcWLwuEZeXD8J5dnM6AtGZMSQE
v51Vn1bereRVni9AVS8OS88RHeQhwawkxwKmR3XmJQ6a4SWz00+0oM8ROudewH0FBbBozgFm5HVw
t2Pdld6qILTYhmm2kqT5r/27EuIqo4sKdVujLSx6bsG9nHpYCTa7MfjKgK+gEqlwSzDsdRZvZW9a
YGrBqbY/V3Ri5WURxDe9tdtS/rmYbnGaTpH9DtHXnOBQqoKIxMDoynd4WHEDuuLDIZsgLo2/GwP/
sQSDmGdTpqjxefEdpibe3SOvJ1oP1FQXW6gk/iR/LszGSV30yX2rQ5mxUVvoX1VhPkdE5oCbRjpi
2LY0OXJyE1tIKSAn7rHWZf9Ttg6NjkfGkpGikHVQXJRAWUzuVEyC+xwQRRx5cHMtcIUjNMowMLSj
DZn5++YGDObjdj5citp0qWn/76UO5wXo0idazz+SIOOWIWUkiJAjdjWDlJA+QFIM7Qn3IcmlPqhg
NLT/7QkxofdYkrX1IEeUAZR9bQnyMsTK6ieqNdxI9M47LwXBnR9++zyWwVTOkVed8/LQagj6+4wv
xjgLNaSeS2MulNnNbWgEYHI+Ttnl5psQwFZWb+jE5YXuBhrf2nSewc+cJwmYkBNhQFzl9hfytx8t
UGxcZ6qD1X+bQc1dnXO975nUTeA+vS2o691P/w9Tp2QDdqVNvGMR7L/gXQboiMDLwNJhUfVHz99e
21fhUBUMGwk8nBPi/48kzz+yUGIqZmLshSseZJv1E/+GbPFcXzUi6frzDCPpPhMpI0icnvhR/Pse
I4AeX/Xl+PB7F02Q78IqlHqErVLJxBzXHgucORIKWSzbOZzkrqncc6d29EGwC1MaKFDPmZUipk7b
RNgGXOr51nTKrjPecutqaThKEH7Lnai0+Lw4PGZEORkPbTy+YPntb7ACgB9bD5DDA/ZhE68wsQQS
HZKcD0OLFpwl1ES1amrXg9AJUq1hdoj6DMegeQg8fT5SQXennJeTe3hNDYh8dMOq0ommGKvoMvQn
FmHpsZRHGKTQ6WmvjpIjOo7320hOare5ZsI7GTbn7vbBqovRb6y9xjcS8taizzonRSLuQ9fbreqB
NtRCFhMGV58mT6Ra90DguBKKSs1d+07SJLFY7BVqnDVPtgSb4niaRJHY6PXZxVLmU+vaARMdbjy0
d+xfl4fn/VJAsiAjfuXivKyqdsapuy6bwSMWKZ7WeT/NeX7tG2/KE7zjDO0a6EvfK3ZvbPMH0mmO
iuryOUzTL8g/beposS88b/Qnve3CcFvFUTkPSlJOvhbI84E4+hpOov+AoUIf60HBWuOc7bZFiNng
A3wi9BUA2excXsFYw4F314myfgZXq1S93/8jWAOc7xIaWfRO0QAhk/Bj8W/lUTkSPcp042fA5vXt
s7zgBFyTXirJTYwY3Tbpsw15M8cxCg/TsSXDWo5T71+QmT4xhIaeo1eIOue8oXfT+64jrnxPzTFb
5wT0roGwnpjIGbE8yAJL4R1G6v5RZwFBxhbBFTi3o3FY0M3Cjqmoewki8NTZ07AYmUNeKj41Cr2m
a2Z5DmS9/0S9IpH2xlU4L0j5WN5pGTD5JbEZTdIXw8SkE8rwI/GrvYJ25Cga1EZPUxn1IGJ4IWUJ
sylHsJlFKJ4oRvk0Tt/525P+VgNDLc/BIH2KtxHivzUP6E/WvAqTL7wjxSUk7Y8Fr4Wg5bMP30RY
G5wz8hSrGQQK5BGUnIBnE5uxV7SuMj/Qwhw+w0pQ+Rcl3aOiPdzpttZnOSSIQPgmYoVU0eSYi8Ae
wAvjiVq8UyKktSSN5vC8es0orChQZKIkDSKI8OBO153lyAXErn306qhbnoOPbJceyh4Q66BXYedE
gBDSf1BmS2xkwTNS9kwyDEK5ShAKi/93wLDIaW4xnWZ2ZzAmgQoNpcHgo9xM36TmZeyVHkz6pgJr
nF3WRyIJLtvU/ICuTpndRXv5Pq3u/jLv9xK3GIda8MhXXFYQtnoVuju49e6lJOMrMYldEyMSZ5Oz
ruiXM3G2SCB1MlULB5JgZGQFN2WMguiQjRO2raGOGjJG0Juz7rHf0e0PxWfwWnOA9faz/NtSRBiC
QmPjb7gLOYOSFAqTfqpVzQsbT1C6zGQCXjNLSyFXMjv3BWJ6ZVzAzwzcCmvhJ1BU3Noxg1bGRE2s
at2oJ7ZkVJuN3YLaXaW76QQlEYjXz3jHSEkdea1Un31KPDku327YeRB4+gWjIP2jYjdKe7HkLonj
q8Ws1HbP6B1pU6j+/pA/+bDKksRj+UHNC1L95F17EmKaXbELkibL6Rdlq6DHQDkCX+KTXCaxO7Y0
9G8Al2nAEUWzTnDFRx6rlV5RRq9EwoefBziI38BUD3z86znnK4i+mN6ItV2ptE5OQELhE2DGn22Z
tGYwncd6zT0TV8Psl+Q3Cw1swLpv4Vx/dpDEvycq4U8KGe2WwZOatNtNKWMYceJSMLjzbvFthI2f
3t2ZQXIQsxMVJTRDobI7r1YvOTfBA+RhRhvPcCHx1idzX9xlv+DwPJHERfsodHx49/ua02VCMGfB
+ECBvFknGDOJ/bKcHZ48+QdJ2LIl3hYgIS5nPUNS9QxFlQljsTAxlhFVs3Hl74e/xSD3JjITwVaY
j4L6uT7T/WOaVZfcVXYQkQoEA9Gz4bwoOsGEhCE0GGkCZZJMUfnzTdqlHK4T67lUCi6iLse/xWSX
69raZ0KCz1AogXTX3q8Lr28qJtY0YKYmWZVaGglEaTnG+eAbqyGhFuEysExK+4AojnAXX6ZrbUTr
3wPM5m46COyIN6LY0SyHnWm9bxRosylh23cYW0NkMDUZCB/mQMDYKX1+b/T0wp5DCZrH9KT8xPTt
pSAZwD0jUyCgTImb54y41m/atuz8mEjpu3UPwYJpnSMIReDcZpCHNzLJ/bUMEvV5WFXqlRwXgrQ7
Ks/NxKQHaw78kIiDbV8dGgSMxE3E6vTJqDxcKVpcVAbVhZyv0E1JVN3YId80pWrFX82PKX6NwgOw
hbCR+9bD96l9yFt8PWThCV/6fnzz52CT7Y98K4dp27BCdx8vuJhzQNz1hFIHm5GURuFwXZyjsG0A
kL6akYWlWkTSXsPdpl1ucGmv6NrBML09Ch15HfqnO8UN8qEQIr2+gzyt/Ve91sITj2GJPP9SUApn
tKZn588Sse7WEk8rqtRJSJv0rRR3U+BTmhNC+713iQb/yoB7ac1PahzJv4t20pwbH3hg5J2982dB
iVo1AoOAiSMoYzggo/EUtwXl1RQORvULAcA5S63a4FmNyHJHK4BSVELr3uQ4ABaD7zdZB/gNlSiq
347KSRqg/cBxl1cczRZBpIortuLSZqn/F0mHcS+v5wOeT36TPGiCPHdOsLNNQzFZ+A5HHUHW3KF9
Jx2tbeLa9jmkjAuu4GVfzVy9QLHXpdvJhqy4fantsFRIDAhDczTfDXvTvhl3oPz9r8v2Xqvsgcyk
W7MFch1A5vUhoKYoNwXEmpScw/GLYMa7Ilkq0jxkdvnWO5OA8ZNMr1ureV+hWG/ErZrzs9SjVjCN
Qy++6cHpHlQheDZLPOPqXsln801SuHO176NqO4YXIYg3RsP/YqqH58y+CDcuY43c2AwCxUKXb1PY
si9x4lFlI+VPHm7vUfKf9xsBUDSNvxMFr5U0hrqLcgWTvzQXXrogvOv67SdHG8T7w0+APQ2UeiN8
Opy+eMicbdIVQXDHBnOeH2Tb4F35j86t1CUlUkzErNr3deRLX/1jPzcPzJUvDiAZu85Y8PvGszOA
+/CHTLBT0MHCAW7ql6kqTe87XjUnluJGzjKXSB2R2HQ4E25mT+q/7RELGdjmeXe8DSVHzTm6wd4r
Iww+tK/p1cZss6ASf3BbT6GvJHDvlCIGnk5xrQUxwomJ12l0cTojKN9swHlXiMEZQU7MYK3ZbzGS
maLvKdxurh+VUws7SWuXU5Buo5HGpuID1kkFbzm3BjeQwm+R+fdpdJfpQNXG1ncTbmdNR2+50WDj
1JbXcENVVLc8kC/TX5JpfBYygyey6sbRGKwNj1NtR71IjgevTx4AxMG0pwekdTsfrEvmJ4CJiNNW
CaXQf+ScfTbgIo3guViTuicJWmXngMf9eyyMM1NzT0uyXOsAKhXxRAjWWrbnTiLTNrNilg32Jjkk
rTgR6OzwT3XPgf8b6JYD06bnh4VI82HwauO8A2keGv5T4o4Rnim9eGfxR+7Y/HE4HKFCn3gG0nd/
9igykQzuDWmxaPqhLce9zKQ/ns8ofU+dQUnSVLG5UQpg4pH2gv53IhTdFUDXsDRhCaM1+rZRlaPG
DzPp/SlwdcHFvMSH6+Ex9fNEybAzqQTKES7jiwRJiMhy5AJKz36HW2Y3oxGEzqPwb9rfScL+IPG9
rWNk0RFw64PIOIU2Dw0Xj+iBjC1qbmBKeE/OrbJxhBdCnnXEVjUuxYa08I3E64Jnj+076HCITJjX
PvOUOwEBVx0nq0C1tVu/j5+3J0siugz/SZu1Lolmdm5K+kgsPRGYv79zO3ZoCaOjI+xFYi2fVwaM
yu2xzYqTmV0LVjmRvXWKn9NbDlR1UriWa48mh44ZVoxnca13DRopTHHQuLjvskYxnaRI5QEnqEuu
P+/kegHVZe37CgCzACp6lRAN/Iq6zwUAYVFqDc0lBaVvF6fboot8DERYYsVTAOwp9zmOjoS6t78d
8XjouHXGU+COSpJ52fVV1y4/3N3lMQRtt8u2GV9kRzKnxqUrmsOCVYo2R/DLJV4/55w7+y0b/iMh
v+tm4f9J3iOfHGygqk+F8qYwHeEECaDwz4UTjcU/qXGxt319h2IR5Z1k4QMycUqMkSF0Rk7b7F0i
I2CZxIFRX0tHkLom2DRqxABGAQfVRIRrZ256QXK3XpVEDlUEPLeyARbYc8HgLF+0K1+HD2RwJdBi
1gY30jPqZIkGfc8DmAD0MwTT+CNgt2NTO6I9oNo3V+3fHsU0YqdnOLQVmS910XVSjo+79ib1khxf
mQKbRAX1zGFKKVOWPUG06mu2GWnbGEOSDK+1RLtbGbO6f0SETidPjOAkpZWTePli6McBKFq7WLX+
OQg55+5aQxRg6jqVackwFRMz9mSH+jPXHcKksJ0rH5yZ2wRiovU9qtWVPZoO1M6joZF31+qUG33H
3f9UrUKgiuKTRu64FfXvOXHXRnS9ozexIMqxa76Exfa7canTVJ6a5Tv3MhEeF4XJxTcZelk1OZbK
Zgmq4QmKHyNL3mfkvhL6dug8dYV72nGHhIY9JcfJpFbySz4C+RFDfa31K3cpfCOG8g8YodOWgp9M
iHnnoZCKOwJU3CtCLxOP0u2x/PTwmNSbEjg/HadVUEF5h1tSoqH2N4t+nNRcGHB0TSrv9gOrX9lD
qirdiS9Q2FGMuBVXDFeFiIp981Y91AJa4Olc5MAEEpc6H64hIIn4brBe0iSMup1u6gQCUyQofh4u
4TXlaAq4BTMG0f52VevAjVLzEdnkaQvmgPrnSBqaKPEE5A50KolGabIH/TFdG9fQ20e2KqMhPn29
2A4JQgElFy9dvb72p6TMfDzHoqu2A3uhHPUgpoyWh6QNxJ0JYg2SFfaY1L+b+KSTmVrOHbnb0VoX
EPS0cQLqNIfbeRdlS5JOy9NeLS9qFizQTwbwXM/Y2r1NrzxSxdA8CUPI7eL8PjEH77cayA1KYzXC
QIXHhdSplAFLoJ8/7JT9MU9i60Q9qdeaxqkD87q/XfliK7vxedpDwZqiASnA+D6EysoBSBUxeLWg
2GbuVPauxo0IVMQp3jo7FnAqrXkqyAtF85mxc+1mQMqchddG+FIhiDr64oYvAv4sz4xb4v/rqxIN
OONenb9patqRqqL027U6TkFO3frMgoMkraxWA4+157TfyH+sy99vfF8VBSthxrzwrjzoCtfFY8IA
XpbM8oaRpuYMKGlnQfCopj72ade/ufmoxbxJahfYrmpL/6hSGrsyc+K/n+zmlUzEbIuPu9Nkfcuf
OusCWaWAWgl/RgBAyAh8U7FRrf6E0A7RFRP1K/M0RBsQZTHI7px9pXmLh8qpr9ywC6asgR8Yluzw
zdyC2FBTjvifUeq1gl3a+RmHxTAuMcY3M/N0qQQc3WW8YOarfBgLJtEs/tNq2PJRK6VI85Hj5ltL
cdYkWS1Mi/t1heXZ/EjkJqyF7rDdLJS1Q3oklkx9eF3amj6mK/9hm8sRNW3wZy2n9MdOXscFJizy
5TCGeFVLxrGwBqk3kxWlKQlpTTmBOEDgPuP3yhCjKdX0qOfEfXgcsW4br0EdG6+BBwoXkztfBNwS
4/aZt/RY8jC/U0WBj865fGYWN7vSLeZLxFiBK+n2XgKgQUShwIpYs8N3ZYBy9tZmwmK6XVmmJAAt
3KwpKIUkO9uxY53qqz97O4WoGVaz3zw1AXOO3db/+s7ujJzsm1NyERcLswiw6Gcs9iFL1zHzcCna
jhbJjE1vvwDX8P/95f/jfVij61QNK/gvHJI8zaYrRdjE1cUFCqR56WwOryFfksbSwsL8v/+M+zsb
MXRYg5+s5JwcvS+jCaw8Tjmle4YMTkx/PKRb5gqStoy/Op7lScf6OflbWa0XYkxfnIFKph6I84I3
PVV05f10+f/uoAX1ZUDG4fN/0I/53IrEUcEK9/TvvDdFlg9/G42jdsm6jj9CYL6XE5X7dW6WGrDb
Qyq1etA02xrn+EKQMMerqD69y0/vdtuMB+kjBzA+LsvUC2xxzsdQRx8xTFMvhm/p6d+P53sWjk6p
bk2Utj+9bihGOvplkMaTWWVc/FBmIE7tn9JzFSFl9FGaVmyk4OKmq98btHnWeQADw7MW79Eg60nH
5RZOv7j3r9NScseJ4OmjwugoX9gCjZE6rH/Os6Aiykmp80oRKObgYSemzYcGDY3Er0yBRq2kgWje
4sy3cT0H4se//CgxAFgy0apX27k9LJ/ZFsfOzrVBN1brxpW351CcfKVmPBDkB6Gc7bsBqAfztDEz
J7mMji6QXF38iEbGhfLoWrr7J+dRmYr+1zaj+rk7sZY+RUjn2TewuM21/zfnWgPna3uY+U+odVD7
a0ILYZtueDB6LjplPPU2uAjbQ8aKC0a089fdL8uzvJmzo4N1HbkfzVbBUt8smuFirBissLCyAWnO
Qq/4SR/Jf5U8A4aB0w0cqj0HepMvqMil/kNRF+i7kymMyeVQxd8Mvw0AAGDP8GNUWsHkyL+3lQQy
8UfJgFK49vmcu1ggKxE/xIdz9NbnrL+4DkTzUpYh/W06RMOgPqgjUa24eOuQ9h25JiPoGPeA38sG
8kcQGKuc1Dc1VAsKT6sSFWvUZrPbfgv8Ul9iwkwMk45A+MKB09qO3LDi9Dc65YzJjeumCIUGbKnW
9iu9zc1XmBGUGjcDj26HxmD/XDCcLSxJvHhyLLo4yEmRyqSUO6kgls4opXxGq5gYOHZSh7r0yb93
Gmnd/3uA0GrgV50htpdEHGtC2M7P4wiDqmh9oD7rtY0dGqqqQhXb75/bxc/NbUbC9a9b+PV+H+9W
M6g8fyjgj2UDcKkYhcDX3zxtYDhWF6mhGVCSYdq8GWlwYeJeDioMMmp7KkhS3hveQP5olZ4yF0ZG
jeMiL5S8DWiqY8qTJLjoh0fnjmlYNLsH11UrWJWKETbCU3wOPZK71M5491JKIvmjPqAiS6wKxQtR
LSV7laNJWMECAMZVePti3EDuy2gJ5wAGGen3P+fXdcpxBT+M5s7GBMNrNh29fmeDpuSlKuCy12BT
Ex5xwntm0iqXgjaYkiv75OQMjaU8BQAKLN3i8Jjgq/MW5T0n9Ckxf6KkEBlTBN7Mdpr9c7teSpCc
M3bJuyY1emNZRZ7DN6ZyE4mbIeyaXh9ljM8jiLjlO6a1GrnKDA4qnqzvMMuqI7kCG2DQR9n3W0TP
tUkEaU2DLFTETY7KqTAKQ0b6dvUqGFvUYirIJ8vAfgDV67cVZfQmm1BXrGkC0O3PSz40UcnbA3fu
k4Tms8TTsrRkDnn3kdhxXF6h8+RqAh3dXBhOb1RpA7Mu0MZ5OIWaryi24v/9VSNuMoyPtQcLtOgR
XMb7TNRHk3cXAxvoMIZs0mVF88ITqVaw6NRm+uYa3qcz2TkRRhZMRxPaNnErj4/DNHL9zVLyx+VA
ps4l6h1WyR/W3pc0XN1j9NXxe2affAreEkLoqs2n2dRcR8unC6vNdmwOE8jnk9B5D/cjHtZWi4oe
jfeHSmQ0cckxH5YvGVNm6ouGmYfLkf3dw8AQlWs2bpult850zxXfYdfEK0vry9k9Fkbio/Nu5JyW
lkEDvZxI+qug84kOXEWu+HnAexQGrg72Oic8bqd/dEXxts0Os7ND6hsqZsLyfB9uyJgqO+8v5GpW
bitmUEVvYG2sk6gZIdYtriscqzdVYWFNtPlzQc7HohbYKmkZqY+80uk+71cgAj3S/cmsAIazO3D8
iz+QBJyzemFOHEjnmTn1WF6HUOthe8v9Rx1OR6l/i59EkFALqrP5+RtgFG6+kTHoJYF3Y1tMM/H0
4ZzYohlzRT5/fpMrZWng2yM5McIacHGTV+/LUcdOmfRf+tabfJYjxVkLcJdQUxJbCGELR6QisAZd
fVL2X5CQFgwIznc32IQ3mWL8nRcTRfdl950vhVOt8lAU41Xvsl7jphsjGWWg0191bYiKdwbtQBWe
utgiOkU03WEsFqyWeUikTKrRND/d0sn73aVwiXXpwOZNBSO0v7DILd2bKIPEye22k8B5buMp+ZDb
K5Qfi51kzu3rlt8Nmg0glWudybMg/3JPS0ygyG+f41xkoRGAjOtmjWL77QhBx9lefHu1rCV2aRwZ
MSjT6aorU9LKNZBnJBWiYXv7diBzOcAwYUJb3BmG/fnhAYsarJ7mLmClbIt2rtSwQTPYPNDD4LZN
MHqmhKe/fbIGiy5bDuF9CAaM44WOhKNJMwrNu5h3r980+q4n4psMJrm1oIsJVHLVVXPwUW4HYgFn
Wm5J1viTyRIe8lkhGpRrEyZ0mljGSyNEsis9pOocl+a//zCgcGfQkvOec7LCV8L2tOYztsZCQH8i
23VWAHSGiGBjp5EPewqXq6J2PhHqWTdxbZQlMBTKO4VOdrZeKUlc0dmEgigEmjT5vpaA7PoRCmzZ
JKrjZcLYETbu3R4C8jKRk+hPksS7RPmWT9pGi2GjBSYLqJY9JqhJwWdZrIA2srU27SP3GnU1g0iq
oBJYsv7NRyOjbsxongo70tZJKXJkO308NAd37oTQGxPaurygSK9f22q1zSt0h8uOsOUdsxMqVkoE
5/gi+triX7VIHjLYtlLaCfolyP8oPMK7ZdftdqUSC9UHO4WCO2rTtihsNjqy9ABPwnQW7owhC4hy
0Ia1+rKm1dQ5RmpkiS8kBQqKFC9gIwyXtA1YS2XTNybvo8Pp27gzm7YL8ofAy7NFl7oaKtoTqwZN
oJNAQiJxTY0MAqOB2GUX298RfnsY1oLMYmDAE4cx94Eao3gmRBrKoKKdGAR3lT3WcLPNG8ytxUDw
HD/5lVHPgPkyhZJR0mLSX+YyiNZHVKiSQ3h/pIMyOXmN9yFEfVZrgBkIFnr0XlWlfc8fKLoa3rxC
btU75yiHUlnuCxXzjydQHi/LVBhcEGP0Lic0FrBXvTZZVFPD8MnShKGNChLvLSFh0/L7Mh94OO64
j4XweFUj5DZZXQ1FDhOCaDqdoqrqOwqJ51kdHC8Wihrk6HvSUb+zT1o3TI5HAfdQnq9sUm2uE3Ts
vFZnm65XxQMTZqHrXAS48B3KGMuMwH4aMWgDkxvBlRhZlX1r92zCZRzu9CFsxiTh7O7rODDtO2pj
dv/snrKJ6ZXG6FhM/F8ynf7GyzhYp0yvHKYR/cZfpOSk/RNoXV+q3BRaNxIxUqnvv94xVGZZqiyX
o01w7H+OiNelpyixBJo4+5yzAH3pTOeM+rW+SF4IRVXF3CqwaYytC0GKzSB7rBXKXdW+VntYKOTm
MIHo+3VjJgyXzxlnouHoQ6ciT+CrhZTosKoVoV1kvwqvGtOI4XJ391qLIjPUyp7YDGMJ9Q+7ICGB
Q1+y9WLaK6yDPAFXE5Z0clXRUSHtkQpVypQUoU1XXXvwii/MQ0wu3+o2mC/Dw13BeGT2KoUSoM6g
6201zbJ7rwCu8JK3de/FdiAfTFnPbGqjMNQsk8TD1BvG7NV4XG3k4PljyLz4nSSzkDuSEf4lKks5
EALrdaK37BP5+1BP/XE2CG29yJsDMvf3t2QYOiIl8JPRg8v8l+jYFc1cD58TKc1XCtNk1jksWGi9
9nDGeHR/p0X63KEa3LAtDY1IVeVOzs/ZXJC2oIKR3JXiS8Pstc/Jp34tb6+vRh9LnAdGg9uzCy9E
b2YCnfCNG9SuL38OIU0tXw6fireZjfQBHPpfIIVCYV/v4bq9DTxC4UJOXVV0b2yqPhyUp0+VDi5W
qGsEkqaxaBqTvbrkn0rkk3jRxJxoW2JcsEM14tZTp5PhpV4mJ0vz7Adjhj/lM8Vwayu4hbJdxACt
SyoMuej/doibl210X8F/3XauvIsqakY02ouxCkR9jFOEklL59PW5JCdjI6wRJdmj9/AQuYld3++d
apIJX5lC4MvnxYCplvV6Nqb4rr90OyHIDOk6Jllt31fwAaOQCwoRfRSZtG1DvLq/6RH9CfdSG9Jo
e7oH0gfq+IsInTBssZtdq3YHVNhzOR5DIgp6+uQiRsUFRGxeWqwaC0l2O8kOx+Rzv8zwtYQK1hbg
DhIen30LNKY9UDyu6HP0/gmuZE5WoPUgSpX/tYLTiQWtUZ399f46LSQsKkh4sHEXpz5299iytAMk
y7xilXgH1YW4xTe+wywkVPw1bB5g932ZwVqozw+FuPm/uEtVl3vIo48UZAPaelavOFCESFBb/GEL
ZhsZycuzfKEAhhwPX4Misl7IMVEhDlYBDLUt4oTCT3aNpJH9hdY/VYEhpi8bTYDIBiUKrgiWdCoT
3JGR3CPOfOQydoczqr84DcpYKT/ZM72olqqjzWXYlcVqok1B7N4FAKWaWyDm33Kj65Gca0Wi0paJ
UBXla/ZTxJoWweTYunncweJxIn98kfbjM2dquvedy+NohO0Sb+wTRL3eqJvBbvOB1YIf08RURfIC
3p65Cybc+b/groVDsOwHRxNY7OoUnobdiSkyGubJqVRlTG3pCeJ1iNCsqpZgWjrEFf+Inktbx4SK
IouSFLWqjGlH7DZyK6IGlShIMrKKETGiNv57Dc2NsM4CsHLtYdKFBZ/o1HJU5jh0/NewG+LCI/IQ
EGY4gjuzRyW7u929S2hb7Uno9JRw4E+/N3xLdNoidtiwFIO6RGTDIkNgIARD8SlqhPfwbzDRIT9w
AV9ONDNcBaGIBtlB7Ub7hmf+OdiixUEr4qpNk4PfBggiS5PePkcOQERxo8sGFUittp0HP+hLf4/0
v1vXfwmpknuPtUTn17OikR92I7XhXVCJP25ekQmFzjhYwq0f771o0aTvM5oS9nyW33ZpRPCERG8a
FnTUQKPC503HHpzg2CFidRDJvrhnvnVghVzPTIMkNGtDe8gM2/7TVTHN83jEGfQd4LeG429nOOWB
7h+dopEJlulQ4snGtG7g8NUTSuQRTIrlEHddE6HGb+AxHTT58l3HjdS5LQ3k0Fi2loqnpU3wnJrf
DraulbRk9iUI7mpk3tQo7S2SsdlS+rdcOj9XJIhissUkWllS3rC6Zdpq8FksNewzuSFTV233xd1S
7K1QvbxukAPVR96lcoG2tex6rc5eqKl5wWwATycXBBGx/OUHErbQjU1AYGef9VGOHLIxzSRJGQcC
zUVSM566r+pjktqj0AflCldOd2R6QxM1OH+PyqPT5poOCfW7xuItatiUkPsY6lMeoTl8Ffwau7DA
lCprI8vElLg+HS2GZ+KfAtf9e9+rAXXP4KJLkx3bz+hZD573hJ0PjN2PR3FVk9ARtxEtC4OSKdPE
3lzau71BpZeB4RI+wx7y6kul4vPJcKXydp19RifTL5qekLS/oRbm1m0ugSG0wkk05AX4Wx6wQMyX
aHtav9FSmx7ZJYT8Z3E+mCFrzQlXdzBOsbzdD/fn2W9BjC3vWkQzx5Pgx8mbhQZFcZh+RiwTovbm
BOnUToN8TnwopoRLp0mvg6xIJHF7ENk23HnbXNRSbE1bfJN2qd0kKmktuCgp3sPG+QFx7szYGmDZ
neQTDA0FoQs0KqUjwrnvg8RwGy2GLKlJrK4Vo2hVUXcCxpr/K5EMqnP7klYLXpDgkCdCnJzqDotW
U6En0OHaBNcVGw3EUHalLldjfDGZUTCtRo5m+6lFHMwlsWyM/XsIUgyXDvAiJLx22nQ5u0ucQwNf
ig+OkWBfANFfWBHIdcsrTxRl5vk9e+Axjmhx/fLO5wvYtyg1pqnj2tSiZfN/Rg6lggjrvCAtIbjS
/VTeKoihZ38DKLgFcU72TA1hoJQfBjra6cHaL/ig4bKvigIAlqPBRd0VtYglf1d0soNGj6YzwcZ9
foI66g+nu1kyritxS8/Uh3RFsqZNw2G3G4aQ4E9xOvS9mo9kviJI4rT45Y20oeO+q9YrIQ/rVb6c
JZK03pAup143NXaGC5g2sUaIWF8t1jYQ5JSx1Y7fPkiRsrurh9Z3+hqcKMp7zlrBJqRUoSwm/sDP
i7loLOiZD430BswQLeooBSNst7dvUzopN4LBWUDXZuanTLOEgMiaWLG+knn1E1UUhzsp6XqRNHqc
I7N+Q8tW71HEfvv5nhtMqp4gYUUjT1yt8LQWpOVBiuF8jzaBRUyHm8o/2skB5QNryM6V0nZkZh5e
r+B3SbPqIpNunCVGH4OMsFjINDczShoQqjCQUBy9ICGEEyYtQDaU6BgbjFJSVQuee4X6GTmZfBgB
gWgftgHnKdYdHy8yZ8jnuLNjJslu9HLDRD7Pt4FK0yY/brmOtrsChnnbfbuSGsmbEBq/d+mJA5SA
ScexGpN1bU2SPtE7kixRB1EOVyWGnRDI3fl0pGb2fAr49ewJXopQlNNQwNtv27O3QhgCAaNT9+a1
Ka7ptQiYGnqAgFroDYd+q90vAgnxJzTl+/TXsSUqt6fAn1CtoE7auZX0qgoxPJjMRfKyl2e2g/35
Hf4buH1LyKHaCQEohJmbb+SXc0AeoYQ4EDtWmy1Y8++KAkJjlz2ArACQt3RPh+DznKoHTKyZVfMw
bKl1GBB1jbETl3j7WJ5A72PqESkflp1Kdyunp6R5FM92HYtZLlPsGEdHCbAuRGS7iePMUQmOm52Z
Dp7TysVrrF8/fHncoMvPkyMDo6c2ICs5jRN3fhXbmQvXvhnZF0+1QfPAuU27wjQ7iL71UcJoXTcD
Pz3TxHj2b3tT7p/xhmJPF+WKwCu9VYQQ4jnUztAhoGKpgyzfhfmRgt+BpaVHsePlFKQbTz6z43C+
tuKBF2qqNPzd73fBrQ7+Z2BmYM6I39q/zpa8sZJ96+5uQAP6mKN1OZJ1NASexkgsqYRjn7HFRqvD
Gb4nwf+h+20SRPTvfONMCeUGQJnzufkANUwtxSDzoFLuOSJPtu7+pnFp7Q8wGSEa2NqmM5L07wx6
ZgmoE2Del2S/Etn2bAoBK1LylSCg+3s//uFNrJLeFGeMcoU+4BCTUgb+/1ZD0KtiYSydAwn7YMUX
VAzOQUpHztFmq9gD5O5EQ+72ozoM8Gs8BVxOTHt51ntXkNRrhNjuK9LkCIDalfhBYsgwTZGYhso0
SdU7L5uht4UfWGO8RxUDhfPsQpHZwMEkPQu/aBp/VwfBz73KozPj5nbm+dlE9e8GECMjZGP/pMJG
ltIY4P/ediLad21HkLEpgoYS08lj8Hy4/tEnkQR7ZkPAtf2OytgE7ZVTM4Ej2MFVJ1LJqOYbDnpQ
s0pLhLJlVkN/8I4EHiJhko2KBmvYsoS+z77bTci+MpbsiZ4KFxSAIc9LKf8zVVWCbv7KGuXAD6+G
ThSDKf1QnERCIxzjKgQILUhXAirJqMuP+P9KjL2wTS3fUdxr4UjVYyJ4/UR1mVj+6rD/FRoKsyak
bInuwnzOSa19nY4wXGnb1mgK1z+1sj495gq0Mr1Veg7pbZvXw7/0RLqJeg0YLY4CakIF4yap6FHt
mQM8VcuPdEI79vjq05DWD1n9hC4iTwdofipOrDPz2uh+mVFNHpWqHL5gHAHCeMkj1JMsOF9aZSuJ
pB6T8qQZ9qSDow3Fb8xc7ornVn6bvEJEvDFWdGPvODaCROA8V0Q4RLq014RbxO3BlSZ0/sKAdvc+
X3DTM9KU/+iC8NB2JUKH4SrITtxUeV95o+MF0n4Q6cnuvtsSSh+BgCU0Q0OKE3dBStUsLn4yp64B
QxVUVkpyYAvPUfIIeSrl+FZzt/PgOUZK0NZFmzQDPguEkgVxO/MFvMUJoC1dmcKUPIdZICLQe1yL
i0mlbvMCFwz08lswKwJCsHU7QhdRckj/eNyC0sjd5wNPqexyzq1PTcQ4BB8pENcgmqJY+5umnuli
I+RGIrR7hmoLQaCWAA7t0+dE7HELXWPWqxgGXnZ9c7UlGjQSCE0JivjeR3ylPSFNayrSPgfTLad4
9jNJ9qQ2iKm3Rud4yaQK2baTPLbjzmNPJlGgsty+56ipxrrqT0H+N9uwtj9AcLvNxn8/OSODGuxP
7KmgmN6I23WI93a6tEAthtis7mVBTf/XA2kUbPMptY8/xUlzu1V5L1rOGHbr4UwC5RJVn7p4fY0K
RHy2lJAv/2QGdhxEQiOLL6C4iAJWXaUfVg9TF4At9uyV5Mg5Fnikrm5tL+HsXt9/piNq2xWrk4rq
LZ2J+9674jJC/il91/vfyfpNaS6vhIyg2bf25RArlZEgHWmrO8kdBIZhR1ImyUYjz9GabNFzFHZ8
J5YAxnKmm3dZ5OKmxqkrCef6YjS0BflX7sXv0GlDNNwkdXk/FQu9MNqi1lf9yWe6yBGyWEKSZUgK
wewj3SbeEEVbuoc1khebzqxeBk4cMcWAgSE5ypWfInNKeAR+o36jbDTGIGjsn66E18Is8/IECTbP
1VFtk3KKb3Icz5wKb9Ju97nh84e9lqMIlcmhG7E7nYPbIOQGqYn3m3iYCUHsZidl+NxbIT5VTmOM
8RPI9tLxx/uDRzYxWUjQLVqqwWpojLI1CHlwtW3hs0w0UNw1PVQUjcb2WpmqRA+uATGV6QB4LFmO
YxphJ+O0yKFvSXdwfom1PgEFi6X0NCNJtw050iUxMg/xci9xVEVKH2W8GOpx02Kn2Lj6+lPA8aY/
viPxnpK4m8HUuYYvd24hNAmIHX149EJzd5OabhWt23T5ZGwR7K+3YH8yE0e4tMmXxJPwhs43TO6K
dCy1owsb0f/gy4CMgLOBi8WfgIbpeqfQUbVWFmSLAwviryCmEGhhKEPq9pvhPozsbMfRZJAiC8j6
2GyyfpgQjUh801cBsu8IMZNYhrJKBLZDn64DtcHLPvbywInvPDD+AK3n6cc/mZitRAme7dIKvfz4
3bhS+vR3ZezerjC23ny6DCbLQqv4tvL8tmE75tDXGw65le8ojhywEP57KvzcZz8wcDJXscUT6AF9
l4iTyUc3PiInGuBUmvfKAZ9Df/6Jvke68XrCNnR140UDEzE6f8FtBn0HDNSSnNZwwg/AplPT/Tny
MnmSVXmvbhCZU6UMUh1yxrSfBnxlDlGSGprdXjbRw8N5FUyQloOc+tCEz8gOdLPNS450qDna+ffV
9VmX+o6Q5o5tlCJDPovBcWbC3Fh0tzcd/lIthyMqiScI9J7/44E/NBduUsjwz07CjpjwoyowuXoV
5oHqyzFq0Sr6vhMD5b32wMIGekS0C2SciRpfdkCOkIlsuv4aD7763SOPHMTjMwhKJ2bAMTnPISJM
NBYdWB4RI1uU9C9pccI50xN0ugTiF3JGPy7d/u+hfJUIJxSfd1+35JRQ41AkUOuWbrT0l8cjFSbS
cAwV650RCkLspDFnCYbQDjmtdepDno9S0fIee6Ee7ufZ99ccVGjZqK9Y2Jygq9aIFvdID6AFL6V1
+5q7fNqvc54GC+/4b58kPo8YIE6CYhwKuQmqi3ZMdpFu6+yQQaiS8JpvKbiUxB/5M6r8+cmM83ZO
deNvaT/X6eTlWWFEjLmuuNmCYakZ1679XW9HMwHBwMose1v9fLVOFGlIB4sje/W5iDPhnTbyzCS3
WVsyrP4TEzBq9N1HEGUvimUdLgsgJxNLfEXAQgHJwubtO1wO0C+Xq4SgeI+Aa8b1YiA2csAlTLMI
7FhU4Gg018OMxWENdWD7Lx7nmwdtGs7bv6FjTdbaAxh7VK3gb15SXLHOlc1OUewdPP/N227Eglvh
gVaPYf+sIZG5PFRcUQw/nTSf49w4crnlbRinYky8ArIMXTDFHolCT2uXfG5irPr3hxBc7mGklzFp
GTzwE2/ZYbnTax50zZggr7k8ZwPWQyOs1PWGrFhpyxDBQa0tA6L1nK9UBqXT7ERkXNQ1BusGY5DV
h8NTM+TyL0sa7pJ3npJgbFUyMVLYRQWD6Uio918P14CLCXc7X3ZOxwtvMzBwjjEbBiwxMyIGWP/a
KGvHX1CcLr489tdZSM2ILv8XFJ47biBMHQPReENk9wXuc36KiN3dKVvEasJaVBrMsRzCVmU3Z2lX
H9r6X4r1Dgsn9oYxatZbzjAEf7UJBrjrZJkew+mTHqPqQo8FyM0aKpIDqecmGxp+BM/oN33EQplg
+wABgy0oD+AAkQok+l1WM9hijEHGTAg2g7qXLv24v1UNOIdQXbGiVclTPsv8w6zhbxRCcdU+om7F
wedwv2wtZaGlATtdNXi7IXAgzbrmEqORXX7m5LJb4H0LFmhAjSd4sAf/e0kcfwcy7J+y7upTXtrq
9yrww1e64vI/pK2IP//u+XisSozEx4kV4XLOTSn4kt7U4lpdxPG93U1O79EKj5iwpSylTzrqjmkE
BE/nTJI4KKiNtQ+yrdUh2xTIrG1sNvhANmCD15kBO+UmLkoM42nEci5n+Are3Nk6Lxsd+H6z/WfD
hw00wy9klHTTIWals6YZlaPisunytQvZj8HYjpPE0qDXVwwUVDqqBYn1kvUwDYe02dAMj/I1rT2B
cezZ3j2E6tQpS6J3Os3uMi50T94MAzLelCxizGJvaDReKmsfVPMFV2BRI6XiQu0BmijQaz3mgZfT
92qbEZDsnfGs3aEhkvspu0wN1B7px+ElFbQNEvbBV4DGPm1HXWEjCeKyDXwJ3aICl9d0xsMLHbf0
HZBeVN60F40zQxBibJkE1I+G2Qbh35M/iMUjeclnnW/sg2sEG++BDrcsTyFIXApRGJ/vZ3eGTrQW
PUG50bGRNoVLX9KCZQ5JMsD5K95tOawbkKJLb711k50qnr/DigQ7FBiHoLV/3Cv6jOeHrTQsSl5w
VqpV8F/MFVcUZZKzoPvNKTiteSjtA0rRMzfwYr1Bf47VFTB4arai/llc4pdd21mmlE16rtF36T1r
Gl5TGF77aNTTVC2vG5u2o+0dpg+GWFT+jivJgq9qN/oK+6j+nj3Cx/9VzlhHI4JtVtulvkOR3KHT
+wIxjLxHdrZvwoZVuMIv0oVpy9Mjh1/oh/dunm6leTsS5XtwTxMC/PWxhkkY5djsrbqIl4vgd5vo
fCqKHOybdcsnXlkJXJxMIeubVtL+Jrn7+ax8monEIR9OxdoROu73hSEz3rbbFOrZP9FpDZ5epDdg
QC++XLnis6IeTg65m4BT1s+iyGb3sN2tM9H0Np9JasgRyF3uTAVh+Q51fFYbBc8oxIKBI3cyJW9+
2+PePKGmXXf4Wg1zjqvy/pAyGAICPVCj0BHbwiN8Zx916PK+xxnpWObUXnEu6bCPBTGSy7H+xLCv
2BIPWwtDcF/+vQ+G5odx4gVistWWml8T6PSUZiSdarMrKW0gIiEHkmQYfF/frvU8lSK85VfUOpkv
Y0xT9f7nSQxOx8BycGUTDFKq0lmGa5vc4sclwSk+iGvgUaH8mLjJleqs7Iva8tZAIRpYys4ohjyr
/Ac3ObrTXc3kMs+j+eJx5RAE9y3KQJLi4+a95lyzqOBeiYdxwMgmn8fsdih8WUhw1oEkHO7B5FRM
6wvyWFBHTFkTkbznTuBJYNxRXZQSbiJ+YIWrkqlBOWNIdsqbT9RPg8SyqEIWBdfu2LajOCVdEstA
u8TR+b9QVrztHO7iCbQVQawfV/cKlw+ZKVJhmHGS5V+PRdpx7EdDNKjZCoTI8pSt3aYjjY8QBalR
8nMzOPIjct1hKPeIoBvtz1G9QDv4vDOx/mneB7EAQtQZ1bA/ogtOfUrHEEPDRRHmjotnlNp05g6u
hCT6d5jsufs9KdKxRumRFJm7V5aXr1SvTUtWze+WDBtByGj07t7E3nrvu/sZ+MWQMT/Jy15uc3Md
gmePIblsRTzDVf+Cid4LJAQj+5OhwuXkOR/1Bnhi2rqf0rYfdkqqsj1gX1MlQj444CM/wk0lNMcv
7pa7vOrf96H2RpGqEBH3pTWdeKrMIjfUNEyGEf49SCVZJRcXSJD1LFVZbjmiOEtb/sKY2N2tPxTU
Rp45vRVwjgG2h2fdvTQB8LhWmGNRVfVGjo3q9HnC9VMFZ+A2UaON5F/WROIcoZTdRkRvTbHAZmBC
6VRYjbwpfpTPTxXCdMlCiO/fks+8zrdk1a99w1NlOJEhpUh/kG/2mmnFbVFFcpsjKva3Yc/J03HS
6uwrNbfVP9Vj89fZOaMIKQuovE5fwoCu/nKkfnSeqC+sln2FuulB80gkKWcAR1QMU66PWXTrgl3t
Jiu4C+O/tBeHU32wp6iSE1YsxrkoSlwvcAJex9s6xrS3pljpzUyeyk6ps6glBaGKZIq+DaJkjYoe
/5be17xjGMaUoZCQGwGRlNrJTRw+Ei5b8UeYSYqA7wIOFqvSaKkns41GGNb47/HGUrKT1ZAs4ijI
uyVkYPirPDM8j1YbXKolCQN9pAFc+n5EECEThgFh5H2NE6JumFY2oybpTYR42EXWWTKE3Np5WrV7
w2A6k7BGjbaeoH0mfLAnYwsMa9g+hmmAXx1/Vhtg9iZDpuNJFIJAuOHWaf3KQI1i9maxRimuCluf
Ni+pNDI17RZMqvZuA1aFvk+hB/JO2+VfpcbCSHTNeLm7wNwmrOcsci1U6WiKdssPhMqijf3b52an
zGRUkAlttFiXKUBE1naWQijIKkYfdn0fwbd7B0tQebnFRLx2opKv3EaIV8O6rS4/i/mx7z8BSsAt
hhvCbgrav0pr9vrcf2YcanMqMCsyEisq8H+hYKPk+92dsbSPe1xFWhvuu8W6mkxqshNwp6nC16PP
iFyduuUV3WsOxHQU6ivO7+1aV5lfjII9shPp/lHKb8tV7N+VwJuO7OSfkjEjjvP3paeE6vcsM7Jc
cXIB3EiC/yELTKoHLDjAtOulWA/2w+lW3jeNGijZuHLEcUD1Iel8H2/eIdTuRJm4rZg8C0SLlPCt
c1smEZGKWjtRJNVwj1sxoDBOiT9IMVgh33vka90k7LbUo3dv1O/GJ+9HKRdcwnco5YlfFkxwJawf
K5YWqNET4cAzNkp6VwLb/ebS0NrSdR4v6wE2xf3uGJVixsvt7J2Qt/dKGyHOpMSq2RVA4dPLmtOd
rI/O6LLH0eCWFsc6sKcZUNLn/nPAmV/N6ynxLJBwCZJCebR+IjeI1S44PK+vOTlW1DJ5NL6K/33y
ltU5XoHtj4whRmvGJKwKBJcmUQyDj8OKrIWNOqlBmT/iEMoBFTk6D79htF98gb9ZmKvt/4ptQ40Z
akNPkM0t++L6wBkxCe9Wwz0S6cUxv3ITywrGJNszJeGNKGFaCMZgiY0a9iWKOr2acCk2fAvjIzJV
Q7tyhm2UFVPMGdRf+4FW5erJDjuVbFj2PbuldhGr6aTcT0yPUa8+BOuGqUwCgOxVmN0AhY9dDe8H
mJ6nvNzVaHvL/HhdI2bblQP5Om0k99gDL+K2kRJylcXQwmSBg6NF0VL8hq8amzfu2AwpGBmSsFAP
Pz8IzrisrqbbdqFTTmhXlVRunzuCi60vpusRugUSViyMuEbu3TrIZFh0ivE2h1tyo20jRIuYxnsp
xZQ+Zt6nM+Rk8ziGsSFlLqSXLwKN+/YbKy8vTC6idIDxW6qanEfo6uVXbZSHF+Hu2h32nq8q0IX3
7ZWGyeN+rjN7fP5PDH9AcbG8f0dIv29Ilj3k3WSAOTbXJmr1OAlLbt+PVUB6O87eupGASDpwkyyk
yMSM8lmimYIsQK1k+bVcVGlRQ75GSDT+D9ONGEoiwN4JTXjw/VYuSRCnbWoPqSGUlqjLDT3jWzf0
6K7Z2ocVLVTQWnPe+mcr4+LGAoRmLFHfzfzoViXIVwh9Uqf3aSP1SsBzUayBTt+OuTgz37smSCqx
U/t4rYixxVgcK6kfmseDYl31+2qmqIuRcg5HXn0pzbwCw2On48gRfE3ZHuZbuQGvj4hh/x/xNN0n
BGg6BwFD1q/vXSrLcd6JQc22UuMFWN3vHQf+sL5Hc4sY+CYTQGr/34mIh3JVw3Tirjapg9Uht5bB
n0QtDZCNbZ1xbQHURlCZY7gWcfsQSoHzghJ6a5QMG6uRbLjjL+L62HBRWhXdWuTXFMOmZnUtQTKy
/vbyTKRGEva5TmaIlHBeRbX68FzYsQQpIQUWI9S4htAcQ1/rWMl/OT2zScngIhViJRyiHNBVwZ4g
uSUQtOzNuEQ8VgC/kSZCu3dHGy6SP8+rmT6lKA2sac53joXp6My9nj2QVVP1iIj03JB/z90HyN3Q
zERq+vFdLUOvj2hWN0m1Q7l8RUsbuhsByHP0nctfGIi5ibem8bMWVJ2lsGGG7ZmUzd5xjTYZS26U
l7AENSPwSlHxBr7HM8Mft4NpRXu4yg0Nc56K4lT9FAgxpThScp+Z2ZGSTC4e1DWO8YKMByeLwo25
BI/pO3JkeT8q6dpprQ7mx8EMQ9KxU6nVpBN9AksmMugSSf519UleUDBMYZNWu2xjvZ6a1f4ykR9L
k6zkhnuoG/C9qy3NJ7w0chr0TL3TNVFA+1nSJ3TPzVpakUShMyez1b6Dfygtf3IzIpANO1tc5+C8
tHUU6drawygfBh5gdN1CEDTDO39PPE278GfF+wMK1ad+SN6f3n+WnqShof6LpUIjfFo6gZhT/eZ8
SNVht7yWgmjkSkCskmzAzlsCg24rYicksSoAeYSxghf7864a9rlKpAXCdNnOgZ39z6o25LfoozGZ
co8fYwIYpsWEGswl5sX6tvzJq/y8Rgm3rWa+nbwLq2LpwgEt8xcwTlTAFx6xZMYwOxMfk7fqZCgW
zugwe+/kev43xm0AcYXVAWE0kBqgPaYHXQZ8686erV8TJ+w0X0Z+JuLtsYCuAdhQYzlSovcsBFc0
+Pbx/+vnN9jpbkq/3lm4xnMC9vXLUkEMSRVJbq/Xx+TD2tJKBEBg+Fg6tqMHwywxaUfH2bzG7tdt
90ZT+IbDVTmb7tBKGY0CBTWFBOyomcppsvZlueFuNV8GxuBvxZ35iy8BOMMmLyilrlV2XAxel3fl
ywLN3JUst+eLlq301GcoszE5tszneAImpoNdMv6IohGi4DVmBWmuQ/mA8w+jbZsjsC0vREsQ8FJ/
m5i8/ASuYCM4REQhEUC0Nad1S4BR4e0y+crYTsSkQjjsMW8OF6+4+XHwCX0YCX0/EtIJ3Qcj13Lh
UfE2VgT2KsPdYWnjP2Lfh9USb01/zBZ8JOJo6BVR7FU5gNfi8VxjEu9EYDS1XEPU/NFstNeGWG/K
F4JeArLed+7c9Hz2tefCSXMHQctYb/cKAaXvBph9uLKKDDsLa9RQSLNjG3eRp0xNtxYe3UX6zAME
BK2rAzW+faGCs0TJLsxfb2IY7XnyFb4s/DC3GNHhsBF60WZQMQHSnIxUJ/cm4YeXYI5ch//IGDr3
Y6HojXirFaYeO2MZE4Y1fn1wceK6S3hFdLpYNFi3SoTkdV5BKeY+X5S6LhpZuyVGvR6qJaA3ecz5
7NhshzifP/MgbVETb+Brpisjx5k8Z8k6qego+Q3CnFb8hELEFwaimlBtDc0GRjaQOYFW71M1WXUs
KZO8PJ7Ix1G+EoW6CVA7qcvIHwRodG8sIX1Bnib47ip2e6wlIp5fkUFXEnsRh/zKywxGLk/ZvC1y
ehXmiEZIdtVWimrQ2xsTMftWdVtmrvIfqffKA9YiqYdyGq4CAE+Fl8KGzOQ0aIyk2X3wyQ1157uM
PRcv1qnsXUrL+Bzs+xXrTi+SriwCWKQLm7dttpIdtQVijKJ5uxGsGEvQzrGyMQfSWjtaCbL2VVaK
WK/E5RTM5tY6zBH6x02xNvZD0t73K8Zz/dhxMbZB2L9qerGoya3cDlniNvunhV1EkmZKEMlc4baH
ig3GQd9VT/AeJBWUpiwRylPuJEyStSwM0FWo8zRuK6lPiKjucpdE/EwPOYAJLg+A2HOvxGz2RHtH
WgBFs2wFEUH+/z6hy0bJYXF3gMhJHc4TIEeJu90fUUOCpXAKrVANX5quUVrUkys+7CNpeS0NJi3x
uYONFBqmyX9zilafPwRsmZ7qVHaFT+gYoPNpHN59PgEK46Aa9+T9qUMLcuLWmjSUt6R3NzG2TOcJ
ckJlNStJb2H78ozKMuZmuutLj0HpdVZhJd/5NOcffBPJxqtkp++P5ppEfkRvPAnwzkKmK1LrsWV6
ZokHCR7cPOkvP0hsqQ2t5Q94aniiFzjPyYpbilvNm1C/Kr762Lu2mRU4mjV6UvGXyzzVxvt1h3za
F1KonY3qxQm7RyQT6znLvzVAl9po/sd5jDQWeJO32OJzfzWm9lkCe+MsM8VSVEIfCjLJ8BVJ7y9i
NwtbNSmiDWyUaXCEUtpx5NV1fcxEf7F+BXTZFB5EoW7/e1uglLK/L1QmNGZQs4/P/MGxIUkGlCxN
nDsIE8v57VdlRyEZpSBXETYObvFyKByWW4a/jsrFH4mQXUDg/UOstaCAKQphODMTKEl+MMF28z2T
+48s8akAIk+SFzUe3BllLnJ/Dyl1CyKY+UFsdKouHvzOPePRkSvq16XL6Nwp/oYYtD1cNfk9gI3V
BIKHXZVI0QXBbAf+9ROJ3B3aXL0qv+Y0SkFuy2HmS9CZEWNHJ8Yydb93N2/aRD7LPajw5yjZBEhg
cGQ5lz0TwZ3XjQrzKQbrVDOp8l5dzEZatPC6eLEnzXX3X9nrDyOBHy7azfj0MyORh4G6TMJY+Nly
o52Lq+LkiewWYEexpd5wGncx3UR5jRUC97mPX34ySLw10LRwDEiQTHhH0P/2twpBofEnb3rYI1t+
8Fr15TrbcG2S2P7U00haoWXDIT7ex9Jnm0YW8wvuqifK01+rLGV0dQTYbHOpJBf8Uexg4pLTWuyG
+h+z8/79r9ZSIayaG/WnzJaY4dv34cLEnEj+Ig/oXTvOZ27pHaVrolV2oZxmmyhTpsVx1BoVbZbW
2H5wWaIkHcAamyoJzH95ITLjwjAsoQYVrLZaZcfXEO6W8+mqpvmHBVRaTfHcLuPDFQkzIRDYH/Yo
MNfUnENbLf6AhhyZxhi7AUOLKlmLXldCG3LUESmeDfTBFp/iJpMj1J7bhG7CLpeSy+KtYPNR1Nut
sJ+rL4WcXrGkysBBX+bRkMdkep/nMCJ0vQTltnIqhLcTxewo56fUqEa9+GiMkSfGyyRWdZQ16PC3
wDEqQDJg1hzJ/18js7w6p809UiC+S8eT6FzWCLa10VngngUcCxZgs7W4cA0lhycUaHLL+5G7nQ93
FcKWHmNvpXEZiGLLtD83osXKKyNq0gpnyFpA5Z9Shw+pdnGgLBw4Qp7VXxUVZXBMJA0w+02dyW+N
TtGZTjnGXOp6E7HoyYFFo82+dCfin6DlMEdQd3kDmm8p/VmImy/UX/zpAB4XWwxKqZ99hOhc/Tiu
dwcuE6wWvTGiIgAn0MHuwHUHgHk1CekojPnYp1uZz/Xf4lcgpjclkqeGapCdDJtpgtFbqCUOJO0k
9icUqLtyPEYtPM+QfMET8YMniIh2GnJqDUEy484Yc1zQJpulL7eZ0LyLUnI1Qj9km+ie0wAn4Iwj
NmZc2JnmAwHimpVhCe/YaimIs+HclW49JTG/0Br6qSWPV8NExxWVFKya/VpdwpFF3rVd69FPssxm
+fe79kWWxpdAVJK0CtVtlRzR56TlDARN+kKznEvjaJf2ddSyQdTBZkWnCw233K7XiOJ1nN7GkXe1
7s8ELe7xdCnZoKedzK0kKwoU8H9tWod2z/BBu/c5WoXKcsbTIVuq4Er3YlhihnJjXP2kRLpcdhgS
2m2PH789xlvJTbGyzGGx6idhnsqeviPjqdcJiepYrKGN6c8vclcvGRzgLMsktg4cDvwHnD7LzXfx
uL59vSjF6xhLVDCT/2aAbShzSHB8I17Skp3zHPBxM5D42SuUefMkY1uHcsxzab92yJDDhiqGdQ+E
//6Cil3Xw6sFrye9quBZzlXPD2PgX8UdQhp+R00ZH+XHq0cQJCgHMzTxjMUyEAeyE7Pf29enUZCU
5RnrJz2OXe9dd6vgcjT9xEYFZXvsLWOhnZ4p7zjqiyRko/FPZZkh6fYAfVwSxnDwv0stpMgStxSM
9mzUJw/vfJI1QCqHq8jJIGAo1m81ApYce9yc1jV6xYX9+7CZYAAXxCJN7C3QSN7UClkXPKUdn/qH
EDYlvLppJXu/GYg8ktVYzaxHC1h3RgDOj8hQx8jsegOLXPoGU9QLrCdvFVGqoeCzvq9AabrGzcJ1
UkZnyYx0+iJ4of4sk2jTjH6VHdQIpe+4THDwill7+Bu4eqxJyo1Db7VREgIdO28b9WYYoKzFlt3D
8hGhdY/xKsHozO8a108Bx4bsyFLbGgbAopDRGkvHyTXt6tbXVmzLo6o1zPXVN8OzOsFn6VDY8tXg
lLH83T3QD6jJKwmauWrXuTeQ0ln1R8VV5WD1VzTfY/SA3RnsDS6m/dRygsHriqweto8YivZiFRR4
NwdFMu4qsSaPEA9hNeULFHWvjjxrTauboW/O3COQhdEziBZkoeuBbdYE14S/HaXkFjKnG1+DiNyR
xyPLNAFjbqJJr6C/BZASPikPXJFLdCB2tEFiejz6XI3BIQORxpLnHJtHb7c+sw8GGFVoNYTIb+D9
vP/N9vmw5H3elJcwba17u0SJnMmFGGICk+DkIpwRjsnrabzTt7ujPp1PdWgocR8Z5Vz2kndae4o2
hJyha8ydpM0BOcySrXi8DDaBZ5wJM4QPP9W5yINT10nDf0l4V96VKH01C/Txo2IIpbYuG5O4xXzs
HJIHuYW112OnPnzqQ3Pv2vII30angI4+L/mBJ1wL1qVuTK7J1FkOMdxTtgnNgz46KoriuFTJw4k7
VRpYYcedM96H9SFB2nMt8qKse0aQOXiiLO7C+MQK1twyxX3SM/ZbdxH/GRmwRemOHM2H2KiZfQDi
t1ApL4XIfuCp9klQt/4CtNuvlx2oP+C64iNlHtBaAYdXXJVUeYiKH6kqVN+9CfDVMARvSjtw6g9F
Xl8hzZwA/rAQGUkn5VC7Tw+N7V+loddQ+smBuMTC7jG9Uo4TQruNKSyqE4KqkTqGZsfDjuh+fJKq
unXAc8jhdf+JcttQ2cl+yzaCstzPfbzAZIjFWc42CEqautFfUsReaiyRVTJ9s55cwtU4YhMmEGH6
GDrT8WT4Mw8jBLP1jlNtPup5z7TnRUpJX5yPnuiHo1JdvybFqEtRci03ISIeFflj/rtIOYd5OhhT
2F5PPYtfTw3aiJm+uWPNFVwYHUf8852LXx5+GsHNRkaT80r2NwqO+hLWBGdNFiARSHZSkjfDANOY
m4oWnzLuEC8gDOuQ3n9gHpcIgDkmYs593k8r/77JpjcFGIXt/Spa1T8+zaEeizkBjEmgjz9yaE9V
p9Iqxvd/Zq66No0b4vB3gqrrv/rdorVRZm4ugwg+TsOi8kumPWKF5CcRhI2konBaVfOMUVbYTQbu
0eyWCV2xtT/T9201QTmoo8sjF0O18IGB4uwchDlHuPYMoSKpVeQNfa2YYxfUFh5hnKjqZweYAt5k
LlRCHZMYR6FnJH8h0z3+KaEB148w7Dp+/i3okithMMvdG3yN/cI2T8rrLa4hcRgI+x0M2NDswl/R
EWJmao0XBGg8bv4yk+9pF9GBeQx3O6c5efBIgnFb1NOB34Si7/a4OjJPfqPB9+er453fnoZ6UXFQ
ppLwlMuAIarJoF/IxOmGWv95WiHjxJkFW7sDnPqeJ3bbrodYkfaITob6t8bx7SW0A9/Kiec/ljwM
68ZDim23CO5xNgWjUA8GdqWGz4Avi9wHMor9vBGN2WGO/r2pUnzzdlBWTrWwVJ2Q9JHWiDpEhNYI
UT6WPrH3x2clMSsSD6cm5zK0+/vGu3Ojdl57bspHb2rOtmYj3k1LqC2mK3RzYRZo6P7xPvLaJHRA
aQ+ACDo6Et7pSx9NuRazzELGdLiDE+sIEw/7z0GFi3BkS3/0OcTZp+nco0otC/PiytwDOGnQbk16
GVjq9XbuPsRuXCEwEfudHU8joMX4vTyhlEzaE6lay7w58tJ+WQTPot/CI51puBI3jSuqBfkXSIa1
ZFuS5ICYF7r4NxfTC0QhVc10q7mGq95tYnW71VQec4nve44w+06fgKRVcR6XOSquyc7EPHd0OAIZ
+D41fAz8R2BLQiAPobRBCsh90OK65LbYxJ9xjRfmAWhlB0wS1s1jfvCuVtSFxEvbfsT8O6BQmIPP
dcSxY5EeGTnHl2qXIN1IoNND5yOWV6mIus7LG/1lxgCNfKnmKyzUhtiO3eVchErqrm6+KjMYihm2
/3ia3C9bU9Uruz2tqHEwapLXJ1tATtybnIQtFt3cP8/yOW5PeMVMyB3iVKQUwBJLDhSfincuteEN
FSVDIGee3o+pLarWADipOYcvRZs3ZCki0CC5+IX10dZdxr+fVZUDbeo5gld8tX14NzVw2N0Tkhqz
ytryz8pBlxfyyE6sF+8IGegmmxad7D+IOYnbF01aLZTjeF9/N8fkf1hIYTrFy925TR1OjPVFhr8I
pHFFwvid748pfMXctPtJ5bXKTNWjHFxfj0Z7ZRlT8Qn+o7FAO5nGcXH/DabMVxBV6fVugTYMsmWo
jdGJR8zvkPDrvIrK3TnjliSYzPb0jkjK3fk7myCYgvjq54HZyI4zClwVLobP1jnAQpP/EtEtyt7q
iRMnzMVxvwodyUKudYpN99Kk5WlMAan3F9CHIOJPAXf2yag8Qzt8cQ74/LHqSi/zSyOT2Y5VdqHf
bmstPAkrF/9FKCCBZu/BRWCMxvPQ3my1TiCv5rpdCKQw50LdZqiAH1ydIt+yrkqg0tzYlqQu4T3O
3BrsqMBJ1TguoJwgS9E3BC2kFyV3bkomMoAjt8Xd/mtbDjMeu4RFbqJkYyDOXURDv+NoyL+4+WIq
6A/WBSbn2bgO3H7srucNor/122edg795FFY0kKidRsVml1HwkxAoPA8Kjo6cCiPcrdAezsIOeSOK
JXEVNpwcjlOkW3grPJGINdLIvOD6e+TETk+sJsf+IwKWyF8HrPxJM2JzQdOanljgpos41+eV2nt2
VzYyTm5zZLhT3Ml1nhieplfFQsBudGo14I3iN41rpAn2iJfJHVyGyE7l978sT43M2fXf0LWjIpyC
jWfx5I/HR8XJaeLlFueOTBS7RyezwizDjgG8Ct8GAvTviRhGLhXbL2rsZpjZelBBb96Tal132sOC
HBDTM1VnfP/07puAbf6NTmp9DunVefcgOJHDuuzULykoaCAz4Y3yUCs0AJOHLW4fTqDCUfGUu5l8
OJEBoje3IgDuqCrE6nePF5Sv104/Ym0Nct99PFT9OChYkkL7ugkmakAQeFdeNjU011/bZZyPXjxT
Lxx2UuZ0aKER/rNqBJB5lhmYN50XRpnvZSrGKjD3a2yP4/YzEUyk7v5vf0Nw/97wpARc+UJIqrw4
UxNTN3438vBatGRzRwlzjJF1cD91tUioE2Wlh24/mnxQrKvC3BPYgiwfsrx99h4sRvPLDgHEiiWH
1fphWAapK4xsDLCAT+MXC8GdjHDhKzhKynb9E351Qd/E/Dkl5rZwUrp92YEsjSErAuhQf/pn594L
oFhnBwFhFMsZU9VmAYE3JlJUA/U7XuLkeMy/3GuTwJULmj2oZEp6ZDdOiYrHF4abXalOUpPOXWn3
x3p9NGIzMWT3bMG9Wsknt/ejLOUPwCcXs90OnHXVFlSK++LMTXEeUnuFHdcNFR0LVkj7wjxyP05l
sJfiwFyx+I+9VqV8u62KqCfp42tjiOsyAd37AoabQDmp7HDDKbA+Mxp2MOYjiefaw7Uvu8K3Cp1w
T8A61BagZKYNQXxCom6gsvuAjcGmJw2XGNuu/QaxPM0b7rrzRfPdkQ+RUiJDl6N7KO/1R0cj2bBe
FC11WfxUMi0m3eqN/GpTWtWEbfjDDpN6G5W4tpQi6fR19ZOgsMMwQpzshFradpQbvv2T8nfgx6XH
ZD8zsC2p+uEPBcIV55e4WrGNBSgeTOAPOUylzKTyrcfwhxvqewo+fqo51sa0S5G2y/Xz1YZMY6/t
lI+Rad2nfQ+xCxpUhY/y3cFh7C9jGxwxD+uhBuJp8aq34cOYRfxoyyriI1yLMgjY5hbp1ObGsPU2
IpjWYQ/DN32RtDjfDc5tS5rzVqkk8vEcdISrSmEQ+f7SrRaCulN2iC3aWtYcA3813PXQoRbanwUP
Q9OqtZm0l6ooVnkqq8yxngue+Gw4uVpdhrwJvmZ2Yg5h640ATSi48jOQriEs+gpFtxRYneISFJjf
bmEFsdNUi8ZsjihZmETQxltAfRRML1R+mqW/nXYC1ECGkesHOzZSTfN8OiNG2H+5eV2P6CCDDbfo
XkIdmh766b3t3DqN16HYaAyyEYLNEOCSK1nUDFLiVT9nQHb4BUByuYDBISPNfheb7rNXeKFSBweP
atH8S6FbGwQS+Lml2f20Gw3xSwmFjCF2Ogq9KSPr8J7xqoYMUP08g90dQemp1v0As6lobrROYAFd
xf8uq5kD0fVjFMzsukCzpSSDtN9D7VoNUQQQz/pH94V5Swe6m3hLZ4NIyt6UNEDkaDbofuVCDDT1
rO3vttNllzWhVu5nZtBYEKxgPIv8r5EFnnm66MWgGmFbOL8Tqt0U5vREymAlhhIs9XHBywzuDKZa
PU4QJTJjUA5ZhGt/71Pk2nwMdiaOMkqV8Kop/5ZWhLu5PC1RBw/X4SAjZW/Zpm/ZzCOHVnXBlrNk
arKd+JabzgXPm+s3Vijv8MLYm2UGSyre1nh2kjs6hWoYo15IHEgsJs/ibtxpDXx8P3Ht1Wb0cQK3
g59fNThHn0iqrxItqlfvlzxZPZmHm/57vMc2VMu0AyWuFCcKAwRSTswi3VhFhv3zghCOPBw6GfYQ
l9zexC7g2KrCl0tKPCcXQARjiqK78lmYH9ynVzQnajG4YnP+6YovZ+lLBfFgR0WyxsMiESRxTt1K
v8yaFpwFZYx9wml1m+rgS880WhCm5EELcq7AW0WJCDvX2x3rj4PCdf67rFK4aNtyFyoKN+LGkVh2
zgg7o5Z748g2llF2/QJZK1MrkyoWoCxb7MfR3IUiV8wpNufer227WFKRPj2tcY2GROTz6RE00AZF
2vw7PWWxmQIAUuFtm8hqcjboSglz1Mm1lrdum8W29ZbphBVZJguoVyVpx/MReCtwppCTjIw5HJA+
V2hGszes1VBFae4odnM3U80U5vTo7fH8YhEj0Pj58iJAQrZ/NGYmLKcZZ+WWslX5VfCKw+9CtvF9
mcP8cgNuUikROrjE41GmDJxrv3PbGbBw0XYglJDKp2QXNOEj/u88UbhA3EJYe615DgNNeOLJSLSh
B1Q85Qru3tgCTiQPvtKKxBmI9cGh3kiXjIxEWS1vLuVwWOXaurUzT/BG9fuyoX+F/qcqlgQ4FOBb
QbcTUZ5Hg1TmFnNdIeWb8mKrd0vEvMG+CoXj1cvUHuBqIVXLrzxY+jsaCxRcRG/cCxkcbmSmZtFS
9UQmhVGWdFfB/P4A0/nPTu+s/zAz6uQEHKO6ebXF7PTVYMO+66U3i/k6FR1/COIbo0T/PRaH/gw3
Utm9VhaNNVlCEzqQ7a3nbThZMqxFPi1ykRL+w8IYnQtpWWeYsEJF+sPJ3um9vXTV6VERdf+1YlT6
yhSltYb08lmJ2TSl51g+T4uJ3Jm/rcQGniwMwyQ1WBUL/V114NyaCMNQt6WJb4iTYQZQa8raVBji
rDcCsWjJ2XmZLRRRY2yHPJjYH1RiuQZjThNrRYVMDn/q9gzZ876uDq6uzDSqooV7qrgZtRSMRjFN
YsO1RWrjF50xo+CScthBkBVlqTzfmbkl4ZYXJ7cQOkVKtsdL8UMceI9T4nnHkeQmmQEZmmo3N1fJ
8LtqGLPqIfh14+wV65cGIvwjlNaWEqRUF06VDG5gW1o5/SjRYk/BbLi8zhG8Ylm0+zbOjLz6qVhz
Xtuv/yOBUUwt49M8CL4kavVuUZluq86x4BPlWgoxwpeTFl2d1p3L2i8u0eXU1cWvKNLHlrrxEgS9
//VLJDFSBZs4wB8hxs1/WeuONXYHOPV2U2bDtjkT++lhYGxXRsI1YRVLm45EVPm5Q5XYLHE4YiPp
dD4zPLAkBsA3EoH4BB1zQVCWu+XBTP/M0e3ACZEbSHbLrUB1+C2+LPhO2EAcen014wcLqPR3zaMw
BJRLL0NVNMsLkmlX9oNYh+ADOENCTREw3P3MY4ok9jY8BdOWvKJss/Oxt1B3Wo7q0IAl0jz/p9Sz
nLh8S98Vm+IT/5zSsOFdns3HWO3ghdc0JiLynfaUwboNhrgJ99fX0AlnmCJXRJA6Iii7G/4mLOFQ
MBMae9s8lB9naow1bBaVD3G4zsn2QFSD/9Fr3HBiZtcXL56ZUaWOGhSYF1NiM5QTWiO4RFWi3Ang
8izmVDmovjqjMZybi0nPUEtLHwPMvGsLXHV9rEwFNBa1YDB0qWa4lHoWwdLOK9EFkUwsnkNcTxCz
4z2gHug413e5VrY9VFRUDVk1BLeJ5kUmY007q4r+9Y0uDjnZNmiRXFlvh9bqk7X5AFv+WjO6jAhh
XHoJX5CJdgfp9Ut7JbYHFG3yWAh69KBZ20U9mcp+0CaKmnuSUijmTdTJ1lUQB5/tM2FlEoJWu7SW
4AtivKAvAErgeHnY6GwAPesdvGYZp7f+YmJdKURHYiLox94BhjJBjTeoxzMj1LWCIN/NvUA1AMDo
wUgKJGDFQzE1q6pGPBareaDw9WXeaghlOlymg9MGeilPk6OVYaqgOz7PJK1bX3VmcNEOtVOsMcL5
ZGM67t2g5vBFfmkmFNuttSFXRbnwga7UlasqmQjejNrUexRs5q3a+CoTgx/yyZnYx0ieW+JnI5tN
AZfDr+NZNK3e2tN5fOrqp3emBzPDMMkmCd7FQJUnQZ3R7rfG2WBiwUKi5f+w9lHYIJYP7/nvrxUy
wX0OkvdkaD1cDcTLuZsyqaVK0yN8+XghZBzQQxgpAtbTciPWOeopZNg5d17chRRHrKsf8YxMWGr7
hfXuINRkmkgeGKaBNT3UOpLVB00wyNXxBOcttFShvcmoQMxDa+KdGGQTIkAbgbtPzmuNSkOMvocI
tCKPCsYFgA0xGcKlNWUOxDI3JBjHKzHQyKlg37L0JHaiNNM1rAy10zEVt1JhOhPxhgG+k5ks84yV
+G63s0NFAHwZxqNebWOC4X9V8g6icAdR8l2h9X4+xvrzK55vcGJ7Q7SADq9JA/uBXfAmmUes0QkR
w6qu+Uag8zSm04lNyDwznRwGqF2Ofg1IE68N68/g0mWhC4wcQWxQs/r/V/iwn/7L1NFoq/MPSnnX
cOX1fJpQ8xsQgPzF0wMy+ty3j/QfRokTFhLJeCHn9cY6KM0zN1KZEWwCVbcJFOXGgkJzM7kXEiLA
m0A1H5VcJpPHULvX1tox/UseRMrUKPI4Il9k1dm4nLuRuvImd5iGs6Cl37UqqqEdhG0b9tCLXs2y
euraheVcNCDe73Htj1WnqnzD2Uqbh+6EPbm9uBqH79vUSgIY45k/JoydpEDim/sPvaUXt4hDzF8D
GDYA4ORHFnvT0qLLrVs/IYDQRyW02WKpGKNQlyEqo7wI3gpB2xuyQHYAr9t19j7DIRivmt9P7Qut
5Ogn/cQeODUnSIxUkJuPyq6/bJVp7K3O+fDWMFI/EfMW0sL7zz990WcFg+9OUMqfmsu8146xW/0m
cg6dG54qTlf2CD3McaYlKgmilbUHg6G2cmn0EKM1tqQkFqGvFgzy2pKhLlzEgDD9HZgcGLqqyDKf
NLOosEk16cjPS5vI3nQavF6I/GXfSCLRRulCu6coJIembs7FUCLsOpAFsmEt3HcNSXL+7uAY7uuo
S3tSX6JnNJKGqvgIbwwuU9AjPxsKqitt9OBgzO0QdOVgsJvSC6S04azfVT/0PQG8zt3oP4IwSPGB
3CvLY0NwVQx9aOM9PdZW/n+6B5kpMrbGcl037XjWYy2LnPEVa7grz1oIW53o0Ol5j+YlOy4cZMhj
U66lblzeGDh+XXP3YvXCdRvEKrbXG3vhOmgLEfQKo2uvXhZ3I8r1EnI92fJCf0bGAep9e7SKlRVz
eqCF6mjdl3BEo/FSh68Bhz1tEF+AZbqWpDp8Tim/PVIeHuvzzHNrhdPzCtz8q2jduoRJEyNKJyrw
M6KYxarDV4fwYUN7i8CcDSTh/+r5tomGXk2vVMlhppebdxFISehNQREJYBsoZOqfz0dNHo8K5VNU
HbhqW6IFr/dtYNVa4IWuXylB48reQGrxXHfd33Q+VAXxsKq9BuAC+Yoe11Z8bF7E1Xtqg6PwCWpb
YsBYiKUdje4O4x0m4ACiLS6f0AcS2Wh2H5BL+IuevKxfwcbib3xzkgTZ3fGhjeYGwEc/ws1+1jwr
r5YXM37nCYsJDpvYjZu7iYeMKgfNt6srHCgzJn8FPC6d2SYEkuW3crEC3veyCURqzUYH42rRMOS6
f5JpZMDGV8RUuALHVhkmK4Z4Hj9HtTLO2f7nxWd0OzrXFyGXatJCTOvzAi7Ci+m1wgx3DkVWQpMf
dL73ilMTwZ43qC8UPwwcvm2zE/L+wc9dd0U6OsXUd2Lx5eb0CDQFjcoe4dSc8sj79NHMt01C7BUD
Zqf3DEYrmVQq6Bq9hmqdxdBQcZ1EWdXZSIWDoiKoKgBFXGyOWfeoyiSu9z72qkycDKj4v5761HVD
9PhS2at/pfA9WZLbs6PWWb+b7fTgkuQIwcSxaMOPwAhxyjSCi777SpMRM9h+HE83cB89gNydu1nO
lBPrj4U81h9aI7+oFSUuAsIYrSryQjU6602phl129aWPRapsP8HpIvLn0u+iFc4Y2EHJhqXd9pjx
+Xo46dqvorK5PuUerLD680c9HLOxv2rE0vNpg5a4YJ85DEjWNsSh6UDFGDZvk71R/pir3DG0yAVq
FHqhyMa8r63EXAuLq7FQT7R0f/CpFu5kBPJiduhtj6oCcnG7kZ2UfGYkERqbrtTKaERL5lPMNqJH
27oUz6UGms3VDigKRS6AodmSSJbgphmUHtnIJHLi+vWHixnJhmYylyqx0iyvVEj2x5H/TpO4XPTT
3RspN1nhxtBsrZ6a1P0dxASQeLumluJf92oB0eH8OZ+Fa9c6OArxiOiSdcaPFG1fFyPibUM2Ry+H
vRbJhya1YnBy9QQRNedG8C3OhKF5p8yTpPJJNsVA6xoTksXT0eUlM35nRDEcHPoVONmF/UmCS0TE
ZfAVV4xaXlA3z1hvCEi9QNMuUlQu7ZG/UAWZPPyRkJLNDSohONIjjpOYgZeQ+a2TZhIRFPNCSzzo
hElscVUpbsQxphf/RGAU/1TROvvoufM2R/QMlTg+jvlJvisyOL+UsHqnAS7G22kNKSW1vQRw3nF4
zhS7XAiDxvrkJl5jzX/Nl2bfBNBhtq26rP+HAsznmVwKG3IPkjRHy3AejHcst1TsW/GIHbcpFV6F
vALlXUktqMvbE2S5isN3oRcZ7/C9alxBsAMDGk2ryf+W0PKIeoNvlKwnvSPw4WLtZB53TDZgFMYN
efcshhKzJ/izqczv66TMyqvo7bfOnBiJ6wBGmnzv5PlfKCKOINff0XzKCc+1cv7MiHX9Uhxrz09u
DzUBKkxzHcRa/hdMModindy0+y92soX5h5xCRAiBm+/vgeG+06qJGXY3bwVqZdlF6NmEx6suxPfB
yYslwiuOvbGU9t2D4XDtQIprq6dCOAmCbskupC9MaJ/kXZORnYH4TQJFGzjNeAVUU5h5rGp0+AWR
P9xXwmFLiLjV0iG8ooJGSxKhSaMpeSrk938sKUSTXaej1DwKLDFp4QYi+O7YK+uqx51BVyLwxXno
Xe4RNmJHyAcGfZs5x/9A8WG5A2ZX9hDVi6uaZzoyAP1ynLGy0nBdC/Yz+4sLhQPXGhLDwYtmmMA1
hd0Bc7Lqrcanyh0jH0geYPObH/dCq/u/gWkDaUHaY1KA6yzEO+mplJFJgi5rpwEEnH+xTi2n3pPo
55AzAo5rLIJ5tZra/cDOQD3EPi/ZjD2GWK+i2xWdwjOKPjavTcbzeHsS+9PGpS9cnbOdzt46Ivcv
9isyoPAL9tMGFejjRcGb8T3O0XOIkemDsdpaaDhhFfY++K7PH7kmCqaE4ZgOpQgSYQR2B6nfrO0Y
3deCyyHqp80sPmhMXVelD50CbWUX9NT4gkyi4PEjvcR0rXV1lBf5rohGyQBaqSiNR4cIKlD1LAxB
6u8krXeKO4BilmKiLO2RjaIMGRt7vw+8iAXMGOryiT5x8VSa3ig577/WPgL+2OuhGx3l/ZZCpuUz
bymZHo1FlDZaY8M35Kspfy5hQwn2CIDuNExeilAIG+uWf3kA5HVQsIsuwClmUq4TIIrAJ0umiabY
lQy7v72zRiNp/3lR212CKZgsjeP2UzZlLiDmtkJ2WthsVhXDmJlQ7D/ZcSZQSgmKg6zme1/HciWF
VPZux0No0qW5tB5kaKMBAGsg15iOOvb7pQydBYpFJKcVCsgOI/sByObdFKXWoHj6lYRR6+231Xog
FPRnz9Q4tSf098Az049Yx+ePkaKiXMDImMyiAVYcjg+pgsVlMQBFo+Z6BzIXKX2QJvhGZ4l4rrtn
Qw8k5eedBq4pK9FInVjFHc6ALKvnkjNmdgiQW28mY7D/hd4E5UBJTIvATyDcIGY4g/2m3mKghBUA
m3F3T+QW7vBDQle0NEKMI/fTFDPZ0sw85nbg+7M5YAUcM6w/SnkPrDniCYgRksoJKUlK7O0vugJP
Ibhxkvbg/1mLTG9bmcdpTHUH0tng/gDmFgRHQZzHzfPncwDR4BKLSQ34Q78zBO4oV/ICHq+T/HQ+
d/4XY8cMYcviueCwT3+7XgYq2dvuhBn/Q4RQKJP8wJwtixLsv4J5ZzNzLktzgfA/wK6nKsvmC5k7
IUOGYW0gPXWAy4/fXDSNvcu/0u6YmrG7HK4Wwh5i315pBOGcPpdrHZ1mss8m/M6DtEmbNZSuqYWN
HUZLuYcF342dxR7sh1TT3+WX2znESKR5POj8JKlx1zsVGMv462segvKpWOaOQ0tcqPaeM96s5Xbz
WxDEafIzUAlZhhd/YyW1VuSzYxdhg49IwVloBVL5tsH6gLCY4HJuhTOYqne7oXJIxUeoAKT0HYeh
0JTadNITEqrqpFrf68oa7RbiJ/mAf9t8BXQ/Qqg/cr9M7FsBLjWgYlhlX4qEDFak9cyJ79hWJbed
+hUd6acW5bU3B72gxyAMlyTxCWySoudi6j8hYUw515ZvpluKDd4PGnkm3hcl5KpXfWRIhUikory9
seMwRK1JTX7HrCx7lyAON1rAtI229+CvX8njXzt9FTsOkXT0oPjbXROvfDp7IcrC7F1E0sF9iHEe
/Snnt9S2MnPoUbFkQ+uGlYmOTuWbIY2/4O3pLI6OONpWCuPsAiw4GTg0+3Coi/cQXCtFdhre5w8u
F7+voZBGGKXB1jpNICBHzTg3QMZuEirniHp+yw7JPPPM8SOur1qznCgPL/xd0hH+MnLWPExcaH1r
SUZZKTQiSxl8zjEpFSSEIOPyqW5+DmOzGZlSXPgFkCWCJQ2AXCyyq6wTeAWU7SVXGaEgVTIA4rPQ
No8gfYsDh2tGN4rAhcDqLwgKESKY1k9DgQ4+SDdIcKl+KsFze08NJpXb/QcmFcjtquGgnfDyl8nF
89M1cQJ9DDWLimimhH5Qd+wXxXN8a6C6MPYiph4M7lsCiIFYPV6yguShBqj18DDOC6giZn4goX29
8s0hLUY4lC0VKvv9PUV4YX+7byhJup6c07cAY2dI+EKjNKOH/1om5YgisFD6v0Dh2Eqhdv8Gp3So
2W9xTnqJ5x8KeFLRMNIik9lhwWH6wAo8AuYFANZw9JwAckDTzZgNgNKBSNW53xj/215rVlWCSGj2
kKPqCFsUX6OzHDQw1MkEO6sL1BYXQosDmePZdeM2iJVSA+Cqswb/oOP/9JN00XGqrwPwAyRjGh8a
4ZU2DMZ3SIaceAQD+jJ7llfRpHe+aDLVyWBQPiyTlsGpsOncvKVHpmw3M97jQCchYXr99ire/MqF
GQ4qKa+pvoamJEsA2ebSp3JN+G0na03fGo/i83Zwqgrn7WeyDKZi/a8u3e0Mi5MJVC3+7fEGSMQH
7gDrArDbSEMOnRBAluiAzhdSVORjwMOyr9A7hJlfqkENFF9tiYuWxAZvkm86vXDJCfHXDpGCKTz/
26cyTrNabVP3Bh5oAiEEDCgbgDSreo0KyodR7wB2XCTEoVhocXW5vBfTadq52eoFbMRI98dAGri/
8UDtYyxUoB7FP7FvSRf2D9gLD6XkTO+5ZVlGlalYWCcimlvgzI7GxhKAbYnuErhSmTnkLwzscBF5
kG7Tg8nS6QH1x7bOetdt0cmuJX/FpifFwC7NZ2iNsPD7VUgN7P+6iDpjskmooKDdeZjjApRvivFR
I0mEJEKrs8NzRpBCxWBwzlTUHfJmk6cjNvQkVe5XcDbL3exjjbWznZmsRnBpDkSxtuS4/l5psAL2
Yo1e+hfqsK1BGeLZQVR8dzfHuRAq4AgCfmrwzKUcFgVjrK7Bx1iY5hcTNKqW+uUfF3PSeId2Kmdm
FLWd8X4ck0OTvhwOK26h6Bu77oRXSElTlkAqwReIJpW67l3f6hACnEeENBmTj5ZpInRzezpgWgCT
Pm3Zt8Sl/foQhtEGj7ceZe70/p2xWv3gQV6zPxz7h60w1sPLddayYht6q2GPZE9vevPNrfjNTa9G
gR2Cu3Qc3urj/COuQDxv1pX7AXNzykHQUO1ZroAa4NcD3Az1vN1rLdh56jEA7cFwxtxmQz7xEpHG
YsQzFe+gjUr/NSKtbv2XKQfdIWI17sbCvkOc1JwArL1FhKA5zII/5FUaO/wD5W/u+qqA2bSVO41A
IwkuIrDjHTDiRq5+vgukPZxTG8TxT1OK0Jlo/4JPpQHHEseYR4Tpr6jCPw4TN3AR0z/6EoGQu/Rn
Tj0sUtCG3/DcWKJO843qpqBdTRn6Y5nLiFJLjdpfPox7nKTjWlAQT8oljW1aMMjHyyYXPK+7aKUg
bfoslYGoWlx4+XXsGCh3gMEdOpduNjTsngODfgLlp1m55AJzbQiFK4jmlylOml/iFJVaHeU23S17
Edus6VXNqt4OgXZWoOrSUsU1xSH7xWVK/m0zXO91ZgkkGZb0BfCkGm3AYGj0HN5doW/Qo6FNkCrz
uUj995WXE+kvvid4GFTpeFIw8OHly3zS/TL05cpGu6gwUvDjrhN2yAShme7bTwUSdX4NSPXDOkOL
zMSLeJQlmyj8ZEjKhQsdyBL5bLdBOdospS7eB+EW/BzMFPt7pMGi3aVfmLrnPAI51j8HnhwWQezR
TyJWZEBJ1MmhwABIHBtnlgMzxpdFMp0V+XbEncsJ384di5vRO53i1ojSPuWV7vAHgF4DfzorDUQw
Fc/y+25yONLktCwL/oYQhx6MLSXwf1ZZ0pf0goTzvDxk5PX9yImIr2WZcf3nZrJ0NAlKTwsBgT+B
LM3JBh+QInoEdu34tfiHssN0utqh15Qb7AKSzwx1ak7NISJjxlGRzGmWpNrjFplZqKc0MAp9+8jT
/AbknQ/ncMVWcG+JOISe54W7oKn48Ji2ct95v7N1nNDFALbs4L2tMJvMyBsGOTSNnId6WBunXG1f
5E3qRd6xW5HjcvKjk1depsW/V2MOUZZxBfxR5bWOOk3HpE8595QZxAE6+gKD6gAs26WwVSQuL36Y
SQJMVK0rS1x2XLPvDPwcJhfzRRUVTR4ZR7EXNzpMXcE+Q330AlT+hs9uWNd7LzwCEPp8aCqb1aO1
7iFcMlhi4QkCB7tvjsdHbHFu2FF8psVWtEGoZuUPKl9P3dqCFIltJvlfYe5YJmleEVpOTUfUI3xF
uYPpbobThKmzo54O9UGedKfpT96GGg/Iw6J+6TcJLF9TvihB6kjJDB8ECY1HIjG+7tUGOCIIEjQl
JKdAAIZOgqiX+kMfq0JvwQy+OHpOUDzF0V9rrAL6vjuRIAozHoovL/WWKtSAa4f4Rs5PIHoftD+n
YXaDId6BOYyfeuqYvCyJzOYgkHagIq5DvBf9vZw6t0llHNHs2gazt+ykZOhO/D+8O7PtKM3HdaoY
sYQ1nWPAdzd8/6TN+6xUfrZ8RypLZfz1vBVlh/a9HNL6y4Tq6f+uHEOXCgG/JZbdV2PDpMlqAXxx
PhsEqBmwG9E8IKIujDaC7XrMUz1soadbpgWF7dmr5tmnQaaTgdV3Xr7zBnhYLPLudjOxc1Al8r13
0R0Ezx4b+8TUn7fB8ageYyrW8nm1xPlLYicTDZjiBdGWU+uz+Agw/yJ+4N6/v68w7G1PMrdJOh/w
69+vS/Jlp2kcryHioH/C/3sFSHwoPeaPEhGDnuziL8PSLZ4azSTnSC85ylbtepI+VltRHpaORK4X
fOFEJpsogLE5DsobYqNisRZoSkFEiJneQQ2pywvbHcr+w9nZhuL247vu8n0R/2IiKyZnc0z43avz
4duW+HcUMRQNAHnTds4dy92MCesQlwQbEVTzm9hQKNzAzOwE5colZS1YgMFPq4zQztDvjUb6ibLS
cNr1DSDODQjiUtofA+9Z+U8PjExcpNSrGO1eHUBrPq7IYW5l6vaboXB8nk/OM4rvF618hrGZj8KZ
5bp4qqnuuvLjcFiPhChVYjK5Irb2hgYh0HtILyRIOq0TOANy4BA4i65bzYchDqwzLV0RrSbSxLXi
/4MFtK4LSczYZM0/Ba8ocTgvQv85E+0eO3VFeq72ZGOAmD0BJRsUraZchLpjYAXNtZ1BFx50NfRN
5trIid2AOuwt/AXoEfIsDBupCSsswg3bZ1j6SAP0K2EVVywX3AoS1lckSE5fs068bIRhTb7yPFmr
BgQNOjMkD0/XoGea6An3H0sS5Z4uA46To/JmfFWGZztHm43Fc8S/2RSqTIjhrZOjbv5rii/QkXgW
FnGRnVaTvZgdIiebJH+kl5aguXx99Hpro3pkPi6DfISR/4qxgWoLhkl2xuNMq/xi3g3BZks+gaQ7
FiVopv8FfaMCHh/7Q3qhOWnWacj048WInHP+PD4FcAo1OzC1buFZTHXyIksNVwNx7Ng3KbCiEWGI
4BYPDqRr1wifyAkjxbgoNII4/LdE1/I/XQ1b4+qQIDh2y7EDmRMA5W5UrIb9KL8XnavJ5MXhJYI4
ztbhL5klwidfyEAsYAa2YpnCF68F0rxcKcbB5Ou4+o+XHR4F+vHydLhqIl73DHfIV8PWkaeGxqu1
WXkTFvDce2TdkwNEqHeehLoBLpU44qaOQGb3I6XAKgh3DBNrTjcLblBnThDN+iaelJ/3Wl6VnXFE
d8UNRsIDDCJnKvNGy72mPuL7x6ZcSMBH/FxdfSel107BWJvlQtKzhjG6X2Inds/YgEyo8Ax38gUY
K+ZBlok2tRxsF3G3PLKkpDqn760K690GyIS1MdQgYs2I6n9IFI8YFK5QgcLRVveYDVDk4RbXlDfk
YG+5+AWw3uUGvkthUDbGzkL8rtRf0dKFlgAjeXSbk4mEWB9Qhdo8dPLbj1keZFO+sLekt+cVO8Fg
+CgfnRBPDcIhL6D4CMYxpY+VwRKJKjV2VL3LL2wHyHlaIIBUKutanEdmRgfQWATyvVeg0vFrUtZM
Hi4oLHftNtIJmY56xYWZdpaDTVRAo00KssIK2CfPAQTEfu/m9qP2OKL3GIa/aXbti8kTiQR3xYzK
P4Aned9G3AhnYaNmJHoXZ0fFIL3qbpsXOWQDEWVDg2BhbPi9dJSh/ZQ1anESmKfiM74zSWTrT6mf
CL282lFOg9a/d219vMNmfIlVQh7fKFD5oZ82o0pEVKqW3dEkpBYrxQ58TW4yPCr3EtaHHf3huzQM
MLI4lE6KQ2OB0HvrBzvse3NVSPG+B+PlTL8vWcB3EWw2iKshcJVjXfS+07sYJl+lkEmOlcShYgeI
mjySBNiragyLePO6SCVWWtJCybAyThqE4jS4n92XNk+E8kDNVz5bvGsrmgTKu4swyT20M3Ao31SW
y+ktlzkLw+tGlw3YIuBV5CXz2Po0mTrR+64DixqOctCIglYwoxDKW+wQ9b7KdXofyfykiY5Nxcrq
DaNo2Fb0fm8Eyu5A6wyPOlF1aBeUih8OBhaG/OWRmC6lXabe1Cn2SknNMeXR2TTqJOTkGTXzah/Q
0uGG8ziGNVk40Rd1hghEkSfCBRD10Ril1YRBF6hQGLO/dUgplJ8v12o5ZW6QXlucg2S7yhPcPVFf
aWrNyC2pbn2honLJFJWv9eCbyKA+BR/d8SnGs6lNXMdOsICqjYFiPEKil9jcuLiiQqXIWT7yLLWj
fDzlUkrtd5eDnNEp2PCzMX7EUbCrshfHeyIrqntZbN7/I8vonlAdbS8VcAaoRf7XXTVuyyyoJeBL
RrhEBKGil9RIYnSOWu2bzab+LdlS3gr71DVu5LfgiAKfOyObVyPTQHT4gKhB4s0bvuAXPe4UusKY
haFWxGgunBdmZHmpe/+akXHuZFDn+n4fnm9CnkBOGfEwgW1qAWEb5mWXzNqBQDjRw1/QuKa1Tew4
EfhXekbM/a3JLxlKj8bRfaojj3mArLu9rUdDud0iuVcfONIgXFLvuZQQxQm+bA+48ZgRfvwGWcjs
OI26saHKWpznH2BY5RdBnGgXlCm1Y6dXUbzAx+hZTVxigcqyTrBDSgPGjXA08EFJGagOu1W7bGts
UPK9COgFgtkPoHmQOFxT3CcEXhkpoq5XllvXO8KRNiAosmOwrm7vtcV3nurzJsQ6Z+CTC63B/oCS
G1zCiw5xtaybn6KuI+N4PI9yqdKLiGqJxfxOIFRUUCVlXv8w7xrVF1K1Z5s0rX/MVz+X57QmToii
6mnt/A6oQD//Bub3BYu77N66cc5haLtZ2GGgL2wG0PC/5i2v6pKPL6OCJHA7H2FTUGevNMMFk8tP
isUX3E5c2SID/HMIpVpzAG0VeCZXiOqJgf/NcE4Rk5Rn6QhcPk124Djl/E3hTaOli+OYXaL0C4M/
dlM2bgVj+2TaULSNDKz6KktYeGNSANfjn9cG+OrVp3b3GwbIB3uZ5rw4YWyd1xz5CdjdifC1zGxa
fonhUr8v0vFwMY2dhznoiUigZqYJHSjUZoEFUqfaebpD8h1fDbqU2/8aGmrNE6dda2KMfmQ8Wldx
vbGF5gpvYWcHbhoBSN8ZWaI9YkaqUzRF9HqwmqBsZSbWxOGjhCDng2lzEaf+K8NMlM8Fw9ppihx5
66LTXxQ5OsSlBVlkDJ20BE8XdFYe/FtIgyd1+4NUEIkDydwt1XnG57OImWqrORctuXsU0r3gMUwN
SkRbqkapbwLLpmU4S5yAd4XTzwFC0L/1uvzFQJKIKk0edu+i1Bn1Bg1xJ8hxAfnBiQUtD63e1syo
AWvcHWF1V6Bdhy1n8M3rnsNPe7fx/d9RCQZ5yCMAPqtmgLOSGGLvcj2Vs20fVwwm1y382rMO0vg7
aNZASL3y2Z6p/7Swci9wscRmW2Mtwez6JYix/vBTWqpBEWk5Cs6+DH4jxsRrJuMxHup8Rf047g8+
YDnpqvqw6DwDoaPdxemUsaHZ8jZvpzA9xUA1Jn9uBstFe8CBYLGhK3c9x853wLE+z/b9bMV3kqHS
MIubFq4iu8mMz5ZXcLIbanghkQ+sBawpX3TgmoCibTiHIvTADwT3IZOpfulThsyP8BadJP9DE405
hkv4439cqAF/tjioySaJNuT7G83ROV9B1+EI8MLIVxVhco5exUi57SiG1X2kpTHNqa8X0GmDT6+k
z9jg2QQD3I5ZuRycP81IWAQIsPXbswMdOWGAGjbr7nZ6DF0d0F+C8ydGBHrCiU9luDLlkwMDGg35
w31hTcuyZ7Q9nlT1DAuUZInGfqvPm3LLHFtJkGrM/S7D9F9CBNNypua5QaxLi3XrNpAwUeh22OXw
ExJOrfE1Md4R1L1Qf5V2RuIMyeeF8BGm/6AoqOCQqcl75eONWugdZRtBGRdSQP8RM1ppCCb5u0EN
rkgrlOczyip7NJ03aA0dvq9b81nP5pDfyENoPyhGCOs43kUaLZ4Gp73FNLn3pzG56nx+ITtugHgs
jQBGQnCnoDWTEVzlkbp/OXFpuD4pOpFXWf2uZSXg1FStJGiBQnxBap62wQmpYMMHdeY6IafWO/rj
lozLhTM2C5tqKyyRITue7alxcrkd4beVwQireF02DhqeFhhBqPo0uwOnOfxKYslsdHPhTAvoIR8w
Ddl9F4c18n2G9J5MeaaBGJ4Tod6W2GY8HIZbp8/gWIqGYivE7x7yDXneDO4TwIbZrE6ToHvGaWbe
I6QxCI2io3AmhV8Etnat8QDJ07E/do6RjTSIitt3EMzAUTL7SN3FH2vOdLs6mrae8VzxPkBVxqi7
LzyzDssTkS+E110AJZcpNgyeWD6Q+WVdDUXa8KZGjhkfXuotjc+LIz5Rsfk0YpqglYwCSMQNrFRa
prgPjA4agx2WInkzFoKPt42LQPZJObYs7FfT99Itn3bV3MO4lUiQZJA+ZVjFI/itG/bTVjWFUqwH
6oByD72jO5UzFzBReSQrqSEf2xmHBa5WqIgi54R6W2P0PgfO2FgkzVnxTMTSc1d2NejMuTxOQEsY
sX+gmK+znAjZLRqWgBrsRnn5lUocwcYWE4eTTrvFND/QjqQDQNdMPpIrhPKaCrUTfZdSTs6erUJ9
2zrLY1+yFjKRqr0QRXsyW9hD2mUB0i62B4du51/2AjuR4nYF+cBud+dyQlALtthihVrTRCHL5lS9
3x4uXx4v7L8q2tdlHVkhIsuP+oQ3Ng5ll5tOhp1Didn1JAu8z+gpVUP0+SzHtWUQ0wBYQ2NUa7oh
a4IyCtpCVvcAVnZmIabMJH2/9/j/YZJyDVCJ8i1588NEjIfEEOjIQcP37w0mbsHsQktbDON5Gvro
D/Ndow+mKO+q40N4S+Ie0AqgoKVXULaqphrRA+CAQxTqIHl6pyoG7u1mEqDQxu+3kvcr5Vk+Epvq
54DWTeEao4QmScmWjQ5ctHwzD8RtZGwQmSuqUVk8sjg0yep3UMPoofZzAFBQhleWKhKy6f4vtmGz
4vIeEd7LASln+pyaKiiBsrVpkJrS4yqen21Q0sbN8k3vxyylCjCcXuiNh4T/pqWlikIy8m1lWeHM
4lV3HLRZwDGxoRHHWCqieguRhotSKgAxHHExCQKbdHHPXlPI8yhDJ/G+uFXvsf2kUjb17xi8RwKo
2a3d0xjTMspahNmzj9RQQLYm2Af4d4jUMoVGuAjCqc9qkDLsNWrPUfELA340f3KDKi2mfl0Lly+k
zGusHsTCH9xGd2RSoIb2U0WeywCy2aw497woDVU4AjxeLMcJ9EGSb8JfKMiQbWbV/T7ErahZIRYf
SWxk5a9obebdzt88Bjw4C5aXjyhL5AGjm0kK8KArmAhh+qjBi/sWDw1ffynIKPGz2QsB/7rzdN38
NlYWgknYOB07a4f+OWrweM3SniOm0pCO7ygW8bQH+jr5V4PxSOhB7BGnFB6Ekkaz+fsG3IYvYj+b
uuN9rTzmlEp7ILmFXmMUz2kolZdjGoqqNrp6uX3Zav3oxm0uWkqdjx/BUN0OS5GMazx9yTdpsOHf
2pUftG4o79Zc6oBPOomtlZsEAUSjhscVQd5suzFWtu+D5BBzj8hKfk1uVgel3d0HOikqDjGvWDe3
uRSWuKqAKdJdjSbebiNl5oYif0BO9HBZyrTSutXGpNkY0jN5RT6L/UZvApAbSrdG8OZadyVa5+UZ
jqto5e9ROH4HcRYPs2ShSRZAQL69WeuAjInZvBJ57VKiNSOoRUWXzloOcC4HoIbmMsB3PjwvpvCm
hziqd5x6imAf7ym9D25bMkCg91w64Zuznlbet/bPov3JLwK8+AY/bkXnBCp30uQ6Ys6qALUR9fiN
nuuylk1bTA0sWvauNVmB8IdWdxd+V82b0YEuPZ0rps2OXyG59m5XhQqQniMJyK5Caiu/jIPutj0h
yVFtOaLp5B3oNkcDj1u/XXzigS90cXPWzsOqvJtshBfo27D5tRDzCI0fpRTVR3xHMCjGtnTDr8xD
7os//FOxkZ/b7a7vMTIp27JJbbJQ/75hY1oKWiOt52rJ8jlzz1c8xfYX7papuQ/udNnGw8sZF7x1
pnNoFtS+xsp7f7Cuo+F+t64vUMLqgBLnsdPHfPUURaF8/ohBxNhccHyFRU38rVUvmgZJGzSW7myH
T8k/8APJjD0pWC09SbuFRjor4zC1dI735TUuzxOFghmY+hLFdQwP6yzrYaCfQItxK7JfFWiPwIxo
YoqAuhwey77/qK0P06EQeYkHCmci8D02jN9TU3ZsjtxhMAZNF1PIS8iqrwdU4sZNC6/tmyarplsY
AA4vofLue9U4Y7VX7vDj3kkEcnrip34v3C9GkcGVsAd9YybK6QgYVjE4e18QQl56/p3uWLyV82I+
Oxatn3upm038QUOBMhFWELv+haI5mUfWKakG37uMA3jeBXwUpXN+o/XGMHni6msYznEdMu8TFsrR
7BEzaxp0u1ycYl7NsibCFvTxXWEeKpNhyM1ZoUT2WSdxMTarQCF/H16j1cOZ8uyRmqJKdwjXokak
6T9XPDB+NPCxjfvBWcQ6ikdW8mTPWRFDva+Z7+f+V9VMjOc4kGcL/Yhqh8o2X07tDU7c1fH5plke
76SFNnNizAuLC3ei/ic/CX/gOnVE7yxvqSOLpod0Cp9be1Znvj6znvBm+5JNWpIcvH6nh9yvBBXO
qO2F0EDcjfeAihaZQy2fCQCvf/NW2PYMdUXdNEav4I0OlfPMs5TrG1U0qbRSMRyetpZEHqBRWBSk
v6sqY1u8jp9Pp/vqyim+xIW+Bu2PujxfG6TUZJKvrNRTGoDbe8HkGJdZWMpzFKagvFrp0cRCHuDa
1RGzmw3jm++tCzuAul9508Gx9yStQ9Ivhu5Vhzo0+4VLBLH7uk3z+OdC/fzzBFJr4sxJ2dB7AaKm
4O56uBHhuoxhePZx/3CjEFKru9ngVFvU3LyHnbxU3y7dgdcmf+x3vg82LCFbtk5M0CDV1ZzL/TCy
LdjFCfV6IPyy1S1urKD2KgH78pYBpN/C/C275pdJlJPy+ZED4uZLL6N+ov6WJ/49skbsX+gEP34W
Qo7BLxaQPo0xXJO5bD6iZ+T00TxEjvP/AFZ1p5a9skBL7CiLYKUHqVLSx4OsxdPstW+BjGpdXg7s
uOECt1Swq8+A7aWEVDvTqxYqQmejsrBWXDQ3P6yCGn+/xNhBJ4tJwFTNRkQ+6/uNq/jWtmNeKtUs
pdew9NcgVHw+AZbbHMK2IcK0DC0YMEov7ScQpgPWfWJ0/YpDN9XrP4xBZ9vv8J0yU7qA3GtFY7rp
g/efylrmT5C1SL5JnruYaCiKxmjK3+YiEdc8jyGd9f/4WvlGUdQeBxpFQ3xJu5WLsYvEWM2peRiB
SOFgvFl/cdDfgE7FVllSdlfeJxNb3iaqUgANjrkEu2ketM6yN89a/ALGjF1GgTBeAoNFpK27N3+n
rN5jPOJuhNuY80HTphtemBhPvD5IRQ7VJngLhXUY+6IzoE1gX9METLKU9Dtc7FOR1CiqWcyuOzfB
gy34lfnFHSfkppQ8FtltCQ8A8bNt9N6sUQYOTnd6u15nW76bSlUTpZx6oE/QsuxgikKVsm86gN6M
ikIEULum3VPoZn6TI/SRtDrNGyN8KjUavzto5vedehz1XMzvFwe3hVZTf5OnDz+GmYMYDWluvNyB
cPrsnAB9KvzQ3LEZGFLDY4tghiRZQKsu79vOAEx2wq+vtNGY//nqbMo/m26+3k6GaGB3bKvhznIP
9jJAe8pAC/0rfmvPubVBx62ELKNKLY3khPjpS19QbdvnWCOTsXa1VscWHTCyubQKPeKYUdnDCpGy
BMWtO34lWyFSIBLh1M1R/DM/7yborW2XgZvwl7SToblzaTwUrtQb9X5zvUFMCwOiKiPEgcisstzc
5UcBw64xD1FV5zCWTxTxpZKHW61rBNJap+A7qe5tAlzv8w5ieltP+gRps4y2p9TpooaVkwt/yhpu
NdXOqeI6rO4U65k3I+0Yen8F7UqkQ77Io+A/J+874KbOPtT8q84U7bYqhvY+05WAWVNpqTJcO+Ry
rwH9jyoYsqmylslHuXGIaRIKgKReasuh9B74ilguyNo/t4Dp3ZgDVte9jyu2cLneDQ4yuqk8L3m8
XOWcTQCAtEia9qND7MNg6+pcsScpe8DEgcqsxKnPmtD0GVErrxr6f1SRHHk9wDtOGIWfi022JQIh
NMRgskblSkpIuOMZHCMs8YKrGextJcqOvqRlCUnW8Ab0rPK4kgl74gKznzldEqgJ3vNVqQhnsfjK
6SasY7VVfyuyqXDfCNOokTGAPpQgQqeeommGki4EjfpUw9ORbIvCtGNYCVOjGyklWNqy9KiRgS/a
nFM0Srtljwu+XeO7SXrelsf7h+QtXnG6WEij/tMlO8Ug1cLJH4xxJdMMkQjU6BiUrS4hKvAzAuhk
McOmucBYCuPZ9U11gcUS3o2+UPxtOjzW9jGuPU3EjD4o0+mqV7msvKgTXMyuwcftdsoIVGepSfiU
CthmJQYD7ZJ/HjxKmN0xM0V8lpajYR2vac/cxxVdW2OrvZUt2MopEE/AplVP9DpQjzfU6GF18QGn
9Or3JeGqVzSGhUBWw4e46itfzBdnpXlUzT3eUtJJuqqnnoYIJfmLHDdq/rBJdDJrByZtLq82C8R2
STgWWJ96ZSQjsOVFsmawuxv3XG2Bks5ZtftD07yxchGZIRaN04EnmJeo6m7jfMS8Wa9EnDpat8Rz
8pSOLK2yAMhj1d3DAbZbnqdXMG8PabJIhBsSq6pPI6A+gbkeuf/wZML9al9hy+pvxxVJB+VAaT0u
lXhhpjFSp1pqoXWme83t21HNgmaZHHf+hw5cHncwNDZqSVXjCDIWuVp9ETH5RjCdGKdoZvgi/lGf
h+eM4XWBjGmadAYWIjmE7ij2i/pb64ev+4V+gcDtzqGkw7zx2HU9hWcpbJrqTqyCMoiKJn2+vC5u
4VOgzjTBqwaxkmTn+gh0GxJ6PgPsOo3Mexev42SSivCKuVme6+VgQTMpqxwpAnbvWGbVsKYVuc8G
B4cU9PxGrO4daMtoAR8Gl0pP1grfPhbD6MIH1gSQnGqklVevDu4xQSQI29LZ/IUYlozHSSNj/kdw
9nYi3z6RgaqYAFICufXs3d6HX9KnOS8nRaiAPmkqN64C1Man2JK/Dt6d05N34GpE26SrRYwDzJ98
DqWxDTkoj/z5roMGLTUx9hRqLmnNc2OtX7nFNDTElcuK2T6r5jSb7+221kLmXDXvvdVCK5LjfJTV
Ow3H/1l9Q90OgmYBA8Z5JUarPlTJ6JlGbBdBlYyerJok/wh4hlhVZO51ehvTgmEMqDJ0jeB8Samq
um/UB+5cetLix7JgnRUQOXSZaWuxciwWkY904WYufJ0DuYGCZXWxFL2ONtWiasTRMsP0d/R+5FrL
lLl6YEoPK5UY1/5mIjQ6knKNIR3RnJlnmH7VC8Ja93rnG2pHLdG+wJLbYy9L1nw+Ift/vk3KY0WS
HthvSnbh2fBgu1knGFq3nEfb6rbBp05qPvi34W58CZ833E0HIqPO4u6vwYstj60wvAp1lQY6NS+G
gjaZlCh0MH7Ti2QgyTCNGu3HdqtEFDk5gnyBxLWUBiZ25SqtJc1WkFJfD2gBms2OnlWzWoKHkBlt
U0e5cXBIVkH/PCt0qrXOlnyKCpo+yfErbD0bw6wxQVqWVK/YuSbL/B4M5pOX8nMkpG4Xv0H3zX0v
OgB1iSw56uRHIYYnYPV91w3ejkMZ21aIdym4DDllPbEWOrgH73QnNxCo3CenVuLYUsm5PQUx13Fq
QvstIY+UHbxii7x9PwYJEJg+Ljx/EsbkDbB8/9DB1kSHdhhsfPAxzYgiwPFObSTTdUnH4+tjqDMo
0r61n7qUgSyfVKsgrMPGCPnlaPyYGB/dy9JCIz7hORsJzLtw2hX9HkOtjRxoCyzVKisVnS5NQmNk
dyyyBxGrrMH7vnBgq2ZGx1AadNFRJyUfn49G7E/2+s5zNZaIWhncDnv0EmoCEsdIu0g/eJRMvDG8
UGVYeSJQ7GuEOORDBTyNyNsy1fKxN9tMXoWqcltIpc3cAeufDFKVDWbD5kHZZ5QPsqnvdhPswhkL
ncGobaGle84MzTO4aVECdZ3J0sRD3/IB7VszmGZP/KtJnYZmjgOn2sdzJjtRDoqvYIMFZ+fQWL67
FH+ghHlRQ3DjEPckd9TEEZvTDvPzxV3mGGdqVSHB4eA0mxB2/iH4Lk8zZGnGF1XGo8QA4uBlh+LD
maj/0cWpeHDJD42MIwcMda9MBpumb3Tw5m2uxfcvPPHyukBJrRnlkDQhuTXZAs27VP7YDDFpRfy5
Zayic/o4b8NEMJC6fdE3k9JQ6ZvA/0GN0vJGwv/yho9zbk2rh9s4uX83MbyJ74rAIsCcM3uQZrdz
fWiujJynhLLGUgOiYCoeCgfVn8oIswZ3O3gr7XoBnk8nIpdC6+EioNotoqx1hKUaGs3mIm8t9jYB
RixJE+Ym2TXDvX5VxMxrDFsb4R1dXPDj2Hr27NxRcvUuOTJSRzHOn0/Z3QoroVLgIJm5rUQZ3rlN
nQK8xb1u8fO7ifRRyvKeGK1sjES1mgg0DF0QmKeX4D2P5l9RvmwHiMCqFyVBShQrU3RpHLkMI7xP
/7XG1yMRdo3pe+xKj1zpOQBycjuvT7GFbbqtIYSzH1DL60l2IMPyZ3ryDoztOI0jcZg5LXymWzXG
ho0aMfqrOahUgtQcRmOLs1vvKr6pTCZoNzivrNxh5Vw4IciSx7BwJ6YssEBLs5u9s3glC30A1wOs
eQmdEUeXnQh7MXvgL1ICxzJ7rs4fMKAmJCUO0nn7c2Rw6TnxGgUf/boM/Hv5sAYtYUaFkrAaLzyk
cVD45TEemuiOqq+i/oMPmlRmszOCHT7FX+qxkZwh3GgEuHMJ0f1xhzRC4u/ej1aLA3q5h7V4RVNq
hI63m5XRRrTb/L9K3r7K2cWViwa5vGG9ofwy3D3NbdZ3hIis4IP5pLdZvasn8iaspQtXrGAKp7V+
Sv7L3zS+20C1Jzh9MGKJNcEN+0CQOtKdsQAm3FboErvQeuxsV5uknfhPuXI3OrkOoIv5NvVzgDd/
GYidSFhBjyuiXRouJm8NM3szjBiEwqzFaFb08rXUfUp/crLk4aPeZUGbO0RxUrn1iVLK+n6TxFFU
vVWe6yx/4z9N3UCdE989oBfTE6jypsHfiz/4xuTxb4GlZoCzEiWvQwtFxA86kPurEsKMnbIV0xW+
spbC0KXR/NVuJgUKJUIFG958D24xmzDJPQRt3AIO2a03eHxb5p/jyIOe4L7v2e5zUhxw9VqbK+uc
dla0aljpkKrGXPQPWp8jsBcuT+aGde815NW8zzFE8ncTLJRDmJUkBLJrHF+swil0y8YiXzj9f3jG
AthAFbiTF/MdE8ELXmofKHTD/k26Jt3nPj763nH3TXQT4rKeV94v3T2A7GdnF6j0vY40UYv22OE1
uVyGvQW63Vl8v0hcArfCny4CThl3Pp2a/j3ED13SgVF7hpAyYqPqgni6AFkVnRSRkEaXcqirf40t
Js3gvXpHkKISSTH9uW8oUxbhHJjfxc17E73XpbSo0YGuAiPhltOLMjZ5vg5W6tTrIxXzVG3C3VIe
UrdFjXhVvgSSz5HPCiZZk7D6ZhVZHlsC9xkar0lqfaQadMI901rYDEM2ycWl9cbwPKSkAhUYy9va
Zh9PRkwYjb4hli37Qte3OCjzHENXMXHJc2ZFPn39StOSi3XI1IVGWrfQc/Nvy9+75qky1Ke3hVLp
XznX13N+VMdMCn9ZD+Jd25xqD1YxV3NQXqv6mCp767qk1sG1kkwBUA4fvOCyTgsvvDGgnKVKnDhx
hB3g4tTAuEXuQRLbx/erXQ3OKwrwmzl47S03MUMzH1cfd9eo2Lvz0a2rwo/x4GSlJH20Lz47CvZM
QXZYPCMJ2PtRosaGeTYmOqmn5lVkYiHuburhyHMvI+aeQ89R4+5GXGiC0g1LA9Z9Ype4fEZPrV4+
gudLrX5lEuhv8Xe5X24MWGlMNwlK9rv7ijcuDHg0t+DXpZOW+VF3VMiQnkCQkjEper24g6hzbsP7
D7N2C7hbN6ppQUpxSd3qjNnSWIpdOR3YOOXIwjdD38e5D72zzv+381sZoq3MPNFbVYbYz3+lvNy4
ZnqtuMnr0bDs5YGIh7HLDjKuhc16GrFJ87MiNsmrYUPZ5oNT5mXd9fWO8lq3EzGy8ceohPS+axpe
0Fo1pYIwQ4en2JqdnNGBRm4vOxBIeTmk6D9qEkCWxW8TUYZWftHFncJEY5akqiDgJ3t3Wb9HVSMI
c4ZIG2mbJhse4yL5h4s7G7XIwxD8e8aqGNj0+WhAX8nz0BqBXgrgcShqYJWof9ZZAH6a9C6oo5Aa
JMtvqRm+aPxkT43xTl0JaC7625KPoE4AwtB3ePrWjWyZnLGIoPUNzWktaRDLnL3eJDxIDqB0Cw3M
wt9wMicOaNOrnKqonV9s0pqsc9+/+7DY1zgdlYd2ujjz2435onwmngbLld7Tmkv3bAzs5IlSxcx2
pMlVCIlh7FyIJygbgMUJ0FK07yQ7/jJLmZsalHJAxQNFmv0NjOzXvUHc4VwexB6YTNZciogN6aB0
GbdUCpQgYNQTrIb2xJro0ngD+wsaZl2HgOpmTMygEl0lRpNWrewjjBYLeiv8/go+O3E6ShiH76Gy
xYPmotKhpysttnar4UWvsUli/y4tWRabaF8NnhfBDEEQL+EcsWe3q3ah8qoqFBWnQyATrRdhwY44
fQ91QW5BmVHuRuuPeCzCA5hf8aZ2rIPN7oyxo0kSWju3nSjzxJ+AOU+3ig82NAf7XqvhzO69JtdZ
4TFQ+vwFpUcklTP5JuSnVMlbnsfp6GSHNVVFOWlqy8fM+FabALT1vZPMqCOyEcOqk33gnyW1Z7dd
MyMsd05n3evbXmi6osqqspD9SMadHwpbmgpNPKshs1VMMo1XimmfvPXCufHrpzwG8haC/55XEsLd
RpwonxRjggHPN+Enef8kfBz4exQoJw/eqKbs84wnraFuv6QQUVXrJlvfMMVATmUgTR6Hn0PHLg+f
3KW0QXyd3Xvf04/UTeKWi/2lF5LgijSta0a2Ze8R9OA9TjUSEcMWXyFn7QWXOBkLw3KJm2ujm6U0
4TvjNmYVyTgztDNy+gCdbW/EdRPFflZlNqWTRPVTmAz1Wz3S707n6EKPI8o2pbmkpFgXZjqo8lYf
6aLAO53o4D2cLNNHrCoYoNTeq6gi0qiRaRB2YWflLXYstISWN0ASvGdAxw3917eCXYoWiGcr3ujz
+jpxVPgOPy1Kz1spDbOW1IBCNUJmEJbSKhoNfKZdWco9uHJQTVL1OCGHidjQ1St1WIqJ5BnO+mLF
f7EjFSHYauYEx5W5B4cV4YuF9+YkOUtVdKt9OVpZCxSppCyrEpniatySBPOL1CecLbQnQSO0TZ7n
Ww4sAO3dSlAKc3yfXkSqPwl6CAyd6Ks1jl6Oxn93Tu68MSXyvjJ08wP2wEeBmfFs2A0pc9T1ituc
ElIXROiF/8OkwfdcCo8G+FTothtgg8lFKbJKEfqayb2sC4iWO39arL/T/rLesVrbK9KxEKn7YcOJ
qSyaKJxSNVVVFthrp9wiErPrjk+AFNEM3fYjtmkVp537A0RKcO/PnBq+a1Zx2Ku+6v8B+6Cd18q2
IxXCS3dYVTrfW1dLsgk1G4rxTC2bHtUqMcUfmgBtaEoCLBX7IkAZYLEQz47675LcPDmCAB2lezqX
j/TY44LVhjmH7yGGEHpcoyfCZs67NFuWJ09/GFXJgufHLt31cb9Lm1ZNPcU8azrqRwcmYFByrv3T
PXCfGsUPmQvwJ/1aJ8ztWY2y2jExnNzXEWUUMPc2qVYLEe4IWIr7mDU04YHXaJq9d5UIQEI50XEU
ycjD9h1YEX/kEZfg0UkZ5OzkntXZ3hr/3/lYLzN/2SQk3bLjCwnH44kgurDi+/1+hPpEB2xyqNjN
U+P6lf/7kjB4LZX9Q/FsOwXGSYjI22DeMTrMoJ+Vml8vaKAHVJIZ0kM+MJBiUL7mnasuEeVA1Y7p
+UAKrdplgAB9h2HdV4o9WtenLXmcaxKiBklNzfzUfJZ1hNfU45kF0UsL31gNlmwTMREdAjrA68s8
Nr5SxYoaDT9B6oWCAjrobcFqFOWRp5F53dDZ75cw5BVhNVMfah95i2yAl+OHxH03uLx1vEP+2znE
umLsebkPFTfqPGKhoOIE1UOez9GP7Q8FJRZt661xjuPCNGqbRsSNDSeeIPPykGXL42MP2svIymW2
Izcrqbyq5QXBKVp9S4itloFRyKQh12bnlcnnw47XazSbT/NTbNQNTBqOTfaYvU4Z5kxqRDnERuHm
0ko/W9Bw9sV4A8tGIM8x8mcHlZzhuY4PEUYoE0AyTgif2ik1yYG9i0wWmmdQz0fIr1g+zU0J6TAq
U8S4FrqPe5Bk4KBorUUb9nIhCN51KRslNZOO5rYxONBYXpMTmvY/ZYc8JoqhQ6xUX1eZizKTSc9m
kxvXIATmDbD1n5zaQhfc2Dm4U+G3hWHg6y5xA2tFvMBv01rhh8WWher3eXi5J3rsU3mQzMjZtD1b
wJ5IyWaRhl5zXdw7Un4im39Dy/Ug0LzF2vlJsZv9XzfaVJU8MgtcVCTOui1YG1FxgXMya20RLqB8
RMUatBGTGzG7UDDOhQ+pR4m4syk8nXBO0WFolPZvgDtj9AdrzvwyGsVZU14hXQZIpQKm6IzuXfB2
e6UpnjrXMs3WlYFuXUN+LniBfocZyGHGzUcYVFZH0F5o1Yz+hOsJjsWCM71vnsNM97lzsWdzqr9M
3Sdots2yDIVJvWx0yIhPyKB/L7MYPm9kbskAFUlFWxUanSP/tAchsapSy2HLM3ghdkUI4uYr9RAP
pf9rvLVHbizzS8coJY45ggZ74ffRhk0WRBgSjCyU7ND1ISpGFVrYIxO6ZcUaS3FaxXVKg9fGVIeF
wjdIU16Hx0GO82lQGCsw8cym0iKJJ1NkX04NJfbF31SKU5h8+Rm19dBxbgR251FYP1B1IcaozZPD
WmLB+uRl4FGIU04ACM11MmdoMjFu+Bug0RWSpv0YVIjEhAVNojlDBmkKRz1MLHUcyntcCn0JCSUj
l7etQ0lGB6Pmf0H4CuhLcFByX4teBjCxf3kF23VAa5gNoQiQcMFy/4ynaCUR83hTmVG0WgL+zXoj
ni0/26cRiiy4xtt05fFMNYlsfucli13ASUJLgqYH2Upxbm7FmNYhebwoxsjq+JJE5zNgXeqlb8ZW
DFXbPWQDHEVQtus3WUNJ0dbAHc6NVV4JvgDSxaPYYe0EOCYminJrzkezR6JV3vawSXyCb2gBMRHZ
FW/58sOFoPnSvUeurZP1zvdubMfZRVtkb5hcAU3fltf0uLZj8l1LvpOmpbz2ylRUIQc7gqb0TXdd
MqTS2SZSI65F2IM2RTNfFIYMrAg8I92E58zsp7rIaM51QotGhMqzV3igdfRs7faahHOx6wd1/aKH
4c6dU2B9OcUUvyFQUsCIhRlHhnc8e3ouLlVB6Qw9d75D+UGe/B5HdOvntL78jlAUFXZGVULFGSbF
JS2H9XN6Q0zGrigE4KbZWKNlMkYuBYaoIz7Gn/ENByWLRzp5M+ma2SIAMJVjKue/az5aH2ocZm2u
CfZW7ndoTKDq0vUu3Bz3S9toXk1f5zOq5MtXCpDs46kfU2jcay4lDqpqAyplimiy4723YxyPtkIP
pF1JkVyf5OuJdfruCQ9rRGgwHJ2UodXQNwRtYlghglmlNnkAZRzfhFqSU2EjabpzPW4leWuzT7zH
Mh+a+gwHcFaFQmAaFhZ5U105LvhNo+h/mKCReQlL5M1H6rvV3NgMmKRmPo/uVixXgujspmFAyvUC
r5H01Y18WbRMeL5l+JGOhyMUp+n3XGl/ATr8VfSjYzC1rnOZP0s6Dq5ch3sSFmkwEZdZoPi0VYL7
C+mtFLlLFp29p29DOcw2nSfNXoszLQFRgxZMnfFnJFrp4poHiGMqmkViOeU33Qp/hy9UtHgh7fYj
IZLig7Ui2DacevUv6R6xGAX5/+sH135cJ7fSZg0L5HZzXE1tPRUUpQrFTDrgiLHEfXm6KGCk0ldA
15wb9xf1jOf4+/vBXG1qfxh0xuz4q59Y4TNZAImOmmLREgIgLG/sXsWyfsSQOIpGZKgea7sxdXem
EEZQUPtO0NcdQfgpq0N0CxSGDqwr1SbSmC/5ByBxU9zzTurYk7wMg7tdfIV0s5Jjn1f7uozc9qcy
9h/HG78HDxIhvUeORgKwJ/dEOg36llAh61NZKok1SzU5VCfn8SJJZfrLl/S13/R22zFlj9pfi7L7
9d5r+lV8DMGHdU6oUbXtJ3BwQI0mPDs07jJ5w6kdn/goghS/scAlpy+VVBdOnfl4lW3MQqOQDnMd
mk2K2tjbEUMiRODg2W4UelCF5/ZUs9sbZB0C6h5XzIGmlQhNhtC0w1KuXTyewmYHr/m9SdjOX3aC
+We5qGJp9L54v7aVLa9cWQ699kPU4c5MzXwz8KA6gbrUXUt/gxNrS13r3fKYTdjFp7f8pzFJUHlT
d+dKGnD57YbFaaZWycC50O0fg28bO5I7QueOWQ+9ApaAV7UleNWWs2p5wM7EI9NsRAaTm/x5z9ox
5vWuatGKdRYH7jwT2zix0HwSTfZKAklXONY47saqFh72gPLUjNob6w6CouZQwQIYKbJ5+PpLaZeU
4U3Ujcn0uSioDs330zviHeKdZUareo9Mr55rAZIf1cLEl+BYhpTE3BWeRMcgdZHGUClqLHzJu8XQ
95OkPyimgFPCf8qQMSC4meVG6GmXZRd4jIKZ4QSt4646ySJVA5PMpP3Mo7VTqDErE0evBWlepuN1
lTJp/He47nlMDkKrp5kkKUcFn00JhO25xw1CCTw36PXtkjyCL3+AYkWoJgix1gpeMGYvhCLOfp3h
hliQ2Dh5L2OJqvFUsghp7GsGsINtMry1z5ik+RQl6izVfrwWmNUBlgu7qZ+VfZqxzb6SfdFxzHkc
wFl3QI61CgEXCswDuPTK3qDad0qAc3bNXgm34cHhUSxpAi321ujWtvXkiFMzx1tZJvtuAUgDriY/
Y9cjU+bh8dhjPekUjgrviGGULFB9dhbMGFzi7ej5f0gubxdM+ym3MheznEJSAUAF4I9Zpu7CZ4T4
ScYYOoAlHXgdhSlHeElragl2L1ZoYFp35sLFd54StcXYio50RuMDFOSadvedZp/vnO7vU9uUbGj6
9vm0vHAC4oAfNVOKLXUShrzZyi1rtJ+ZEsG59gxsYDzrqI326MBDsCFloAbcU03SwobFd7j0Z0A8
LaXBfN6m/6wELBroloAlw/bwPTelpOq+kCUcC6KkNaX5M5g4OF771jGmbuA7thZyRfq9+Rl30clG
y7qp3T4+LCXy8o2FiRX7u2GCkKnkiv2zQEe1zHwtNPzAFcNG/g9LE74Nd4iTdOyhzk0EIW2L1a21
GH7vkPQX20mr15yT4dymBC8uPHWE9VC9SzMkqjFR4zwdgJoG9RroqYUbv1FncQgPESEymHAPXMWI
rjnKY0gBKskoL/2uHKvv+fOXMx9TUylpFHsoKpOEWp4BOTOl/3TChOjGDbO2QwJlMDJBFCW7YPLQ
GuyT9lT1s+zMPU5eh7iU90ASC8j/mzDvE5OfEx6qQ7SKHIipEos7Yw+fFp/KkAPvj065xFa5TVBe
Ha5QLY4zBTQFWY1zCsRj2gO0QstfLAfl+r8UjjccP4DDIfPD4nAn8AkvWnBGIo6keFkDA83uvDFU
CcSvCuNRytrDvnrQ8XjGD/1B+fluhDGJzFzLA/ax2haMj30vI394CcZYKPL80Z25fu7Ourq9+gGF
1glOGObS7jmz1Dq0562XOdCbf9G9EUBAWineZ/e+4g1UbvfdTXP+A+YAoCy/Yr2TeLDv41T+M7XG
Hzc565BgClBjRFqF/MpAw3M6pnZefT/lMwNdBvZicFDTOx4ARggwXSiN2v5a8HeigQRRXL8Hsill
aFPs3NrIooKgc+nAtlECJ7TyaAa18g4FBEnt+GPOk8awqMwUNem0NnEpTOZkK2FZkHoyDDkxifCU
2tRzebgRXNEKAK95VAqb+tkrq+ts2s9/Kks6erXjHWeLERVhitTBgH3zWKQx1i4Sz55Y2+fH92MH
0K0Qs6fDMRY9NyxZUzU5W353uGQfM1RhopAiEnoAhjP1gaMXk1qKI17vFddU/yr1nw9QQOpckOGY
4dyHP/h/aKXgjp6DmH+1cHxIDqO5QDuw6t+pnPHUJxCcvwYmzS/sEZBqOJcBmp9HcfsuisZ5Q7OG
rDpnF6RI0RGRlcBEEE0GJmnLS++eO47IweQsF/b9OXivjGeuAMRD06L4XyhciIeABIOeyzqjd2fY
9nSKM+SuGiXfJO2MYSnZ6xlsiBu7YcU+6QPUouNp1y+ya5tyQUyarg6zkM7gdcgqTSa396MmUkyw
DG9qhlg3PUcnF94Bfl5kNwX25MkyCY/IgODEllDFkj3KdGsOij4KtX8NIbLXXPR07X+S2u6zP9Xa
84c98aYKlBFkBF1y8g0fRD8YB/BryeHSi9GFtxE2vVH15a4Vv2Uef/wSyq5MvupMMvgnOQHEJU2i
VutOGPvT9B48aNxiiD1yfAQSrU1W05IdVK6SMvGsXwEiqCQJqG59ludlDIE+vFFaoiy9O6+Eq9ot
jxco2GEhdG/CUKUSWMFY9VIKN+dizfGsWCGrpFvmpzkSuPIltN/4IJBm8y6UczSlp0PkkEpnj3o4
AyJMi9SfvXoRCxf0tpq+8Q7Ehm6fq9dVY9ZGLA2ZuM/JOMLa1NGc94DT48RcD/GC67Hedt5mDGyU
nXlNEhnsvQJWIcveVTCEU5vuVA67e6qEX+LvRDgeiLG1CKUtCx9tIQTo6AsKClTF0CZRIbId8AAg
lZC8NENO+j6whsNQWRnc/y7AYr7hddGdAszKQe8HUrxuJ0gNIFck9fTklxE/vSwiGKIP7OA89JmE
7cgLlhuCrPJnGTwL3FIKEpLRaLwkCl/nKTOfDAT1HmpLMFvv89hhDx7wdSUiyPnwAhL/7BTHfOxr
edXFQ/JiBzOp/W3042AdGsu1LWYGLTz1/Cm5K4EWe3nbiwiAzW9P+wPWD8S3vo7LYxRHPzmhiTgq
9V7MfnMbHC6tWUEaLhkFPQSNwpVNX99Z4BGvkKUcqwG3FISt2ysJMgJV4PgFOVHdZ+vc6DJlmkF4
/POK6IGQvoas5bheLR1JOzQm/yHHYalw2UjmUTV8Ks66ouss+kjAWuEXtCzKJfjeH8ECTPO5A1tQ
x334V1gij9Ocg0Ms95MaGy0URkpty/JdP28teULomBhIIR1RyBRFZCITFsKjXyx3uKO+3i7DK/bn
aE5/ij9p/lAIAAZfu/WLHMJNdbxHYPhHllcIsTpUa09BpTCNVYhIgnTbq7JcZbm6gpvpdGao1Ed7
gVium7vcAK+0gVBjYZc4X+SLR3ZIf4ZMRzb7veuE2NGfW1IlvHjrbo4820dmZJNR/oxTUuDzGdiL
IC80/HNvhl9Q24Q61IuYy2ct/67jmT2gGmxyIst9jivwRWd6ZW0aFNMEOymu8ViIY90MQKE36ZgB
yt1qBsmAFNXwDB72pvQN4wG1EKgoAnPKwCVVbUQLwklugwPRGQBP9uvqoat73mSbe0wdEEnjB+cV
knsf+J1UHGe8tijM73y+WQvFZ3cD/6Egx1ipaa52A5fdMI8LO3vATrsvOOIoze92JngackC+pn3v
Sxj2l54Mstf/P22x1FUee/OrGyMoV9mnhbJPEgdiDBTN+St8AhmjlHKMzQTcv/9E2IvAoWaiIZ0C
ylhDV9irLldDTSeFYnjlftgnc+Va7SyTlGONKUtWzeCcGew/oQR/om9SGwW2j6mmHW5NirtgoXKA
MZzTPG3P0DXqGsITw44BIb76fPLMt3ie4HbhyDtEtCV41wHIgkjELR7Kh+TN8doau48SnG+PVbvu
Fr1KO7SVBZed5s2F0e6fyzm7auxnE/Ou4iiR6fqTH9sWZJq9PxQtamRmdg4ynoSE32CPjLM357cW
lqLfaAZyA23t4jCXa7khBjwRjhlyRjryIioUNRea0+n0hponkXbaZ42q1E8R9HaYihJQODtEQvDQ
LZaF9fXRq0ySNh7Wtks+a4XCmkwy38Nufc8bCQzpMG77LpwV0bzTHPuiiXQM7B4R3FckQ+g+BPVO
NzRwYume86ahEwpG3dpu9+MYRq+wNptwQk26N0XNQ2gehsMIfAYPH9jSdARIIePuk7G+xt+E2J6p
fWj/OyFarMv5hM9taysJbh2cGbjToB7C3vulZO+18d2qdTWSBMpDaa00etF8mxnB3LI+YveCukwr
Phs8kS16qQ8XOp8gesq0Ip2DPI+il9TLtWhHTFbC5kQmR/0f35+yR9wBCkn9aA55UU48EphZYmxm
t/7i3H35Rwuj3YKwO3G70djh1cXwaqkplhSKHU+whYpJw5RVb6vBE+8NI8JqnpubiNQtu1dUvc+f
7f+pSNaw1QJ6A8H2j0m3dJj2OSGeCJ2P+ACDarsNThgmNbmWCTz5gkPVarWHByor1e8x1BhDb5Iq
O5I7yPdAiKDT559/0dCuQ/D9eQocQQtY5e/ZvUpBB4ISpUIXga5dKwCbN83+2DwZX7oDDX232esm
lp4TEexz5Jl6snWsSXZUtPqrKi4kVasN/W4Vf0GLl3WsnJINxQxXqEMpujd6ABgybwdjrS3tAFa0
p0YnD2Dpi0HTphK8vNDXvAGGwq/wIY/veB6xd9y/y6kS2aqePqK9HoHdt91glmBWB09DHT+ppnXH
D8GAuHm2eJz1lUhheY/upyxA/dVC6HfFZ1MwEp9lgN0KaMyNH4x2sUZEnGY9IZ1UHS9qWlciIaod
QNwR88eDvEvjFh4EoQnAW3UzG0a1r4Y1JJfGE2DQlWRRwI1pGnzSq1mWmg/ElWY280PRIDyS97oZ
fiCGzyIaVBnDDaSZUjhVJDOiz5EzyBWlVdzCsGbvHdO3qHEa4VbTdu2DZb6Fv7+Orf9ANh/NI2nR
oLAEzyz5XIuXU8A8PvgGd4xdTfLfjj4DmfyfnxE/zd64eEfeLqTsxX+4RimewOkBgW9Yh88eJ2yV
jTk6nRabB6wnjmL02M769bo8/MmuB//+ca4MDlwo0s4A35pJeF1YLjeLJvaH2vAPjod6dM5gUiCY
h2JPobCjY+2SP+zxoApvmyw2qNBStaCISX40igZIEEoxaOFUJ/u/9oauphpIyplJNVaCrMDgyi8+
KwvOzskJlzP9QVafRMU0CZBIWyyWjqmRXlFVrJdkNa08nYlXIo12MFwYoB1dnbZXCWKGvPs8B9Z1
5NSSQR/ej5T5aGsHcaxyq26XQpbssAiAMPLpmIn9xvOXIZ2kgf5G7syqDHi3otwsCLc9KZlB0P36
ipWWpXTxSL1TJcKwp7Fzp8W5/DQG3ucAVAyHIY1hNhvagaPPeoIh3MX2nDrCtRi/XqbdW9D74LHW
hE4v8M6j1GuSqkiuZ6wd2qBkJ1WGT40dEU7GSZr8vZAp5J6zPUP46HKo2Da2ZrDZXrDxKRQz7X9+
yCBoPAO4x1+0v3JzUef3jR8hTX3KgCltD6qYucUx9ygwiCnQ3hw79fTlInv1nkvekzh+U+sohUFX
Z+4MkOGlGqMawdkyNYkLph5j1rVjpzvUWp8Nqzwp24cUS6gS1hbjjEbgj6J9uhKMCsgu2AeWe/B8
jY9Qllfrs30y7sElyiPr7tM+t02jduzGKkXpm5hFOhglblMaj9ICTh1Dg5z8Q3YXSRnKb5Gt59lT
eT4Qvl/CesQ10zfxqGmYCR+MRt7mRYwVYT4oyILou1zXDU/juwurX5Yko7NjCPcKJXVrIV1phdsF
W26n0PJGvZcX5EUSS7E9FwUgXz/V2Kntoj4BnXYFmBufZ8XlFxNaVblasHTHn8j6pFpHMZUd0aAM
q4zH9h0pWbAI5l0Vhumu1ZUozUtkU6AoVpVZacIWdRhuAVPkjnXs7f02dY6+MHdnW/SYFBTv27oz
KSG7pk9VDbSqMC0OxLIgtjeHztSo29yyr1uns5xNGealYZ0bQ8Jk/dGVnVIg3724Fd+fRFoI9D6F
TMYOiJTs1TbZR+gweO+xeobQKMzjKDWZyprL9nJ7gVdFvAfKRMC7MC6HqbuxvpNWbnltOQqbfk/o
sJXFdrw+/wUz2ngoQ+liRXtp183q8+ZXu/JE4FqSJz4rgEGiuUbpWYN9y7BMtIdV4mTpzq9BzHBT
5pAz4RITs7uuiWVDND9n4CNNJ/u3qQJCMStcJgHpyFqt/gcWDIiLc8CpC9Jm6MfjGa2K5v9RM9RQ
F7MgufaJtDuuO0xxeBCFPlhXNmQnYi84I5SndeQDr8rJuA+B6Q6U0wlo8McCTKYEMkJw6Pc/yHmx
QJF3XLpfFBRTraS4vby5sjMppqK87c0oC+GhiZo1kuvSG2NTXx2PgvvylbVmsOBhqvwWlbr9LiGT
/Oc9pa4iDye6JmJkoJ5ZoFAk+hV1+Nn1gKYZnGXfHOC/xbfhYZX/7i3NDEsqoPUt7nVMZ7RPwXko
jYPhbtB5BUHpVyh/DQ5Eo19UParMVg5Ux7zE/njnZ7FGkxGl/cCEXRYZqd+sd1Gpx+HJaX/OxIY7
C2EmfROxvf0HX6DyEaQ2fEHV+JE7cmoIzBHSHplAKKnZ+UBidk8500EJpHSxrn5FdrDlkdabtG22
GxT/P+loG3LtVwLrtiMfTiiDEcdnRt9YuuMuuRwMslK6rDWHcr+czUZF94VsfSBRL9pVW+Ajox20
VXPiG4vlZ7/bSDFrvjz4OL/HKUKt73xN4g8aLma3ZpfHazDgnxNDkk/Ueb5lQfQr6sKLR/XqS/ng
PLa1Sr+XA9i0yQEXYTN9SvcuzbNjhKDh0yGmMTKJHe2ZX6xLBX0Y3dbGpfrj10rut9T0DycY2jlJ
cPiq20/vQQfeo6Uzp/yfBg6yFuiINnxsxvyZVDOVHXIgkcgxAs3kABLUip1eiQ4NCyrKZzGikdPy
lScqDqE7S+dhOVrnf3JoxrAKTKgX6u9cOXTUt07IEu9fDDV2AqG4TCBlHNb51XDDkx08WQT+0yxv
slIFDIwdz+8RB7kJxuLaKVhJP6WGGLvDlbpktP37mDYhGs2ACB31CG4Sd1F1jJYuXMNEgq3KgDQw
LEFVvsa4+rVsLUuYbrQRLuPPsbuqWDVbGOOHdk7VrS3OElW3F2U45R8J+Um193PIt5bBipSvfMBZ
veLJ6L56jF14UvSggSqLl0qihsBKk26RoKmh3fYd3bNAJwL66NkBF2y6dOgEpu7003rqUOyvl043
XsbSbora07xxCDTpzUsh/D/aP8a1+uiPYLCR3Oy6FNXoL134vqAZC+f94KcSIEuTu9hR3FbrQvbF
A5ywkKczQwqruFR6dc+dkCeQTObZaanJI2Z5MZ+IPfWkaiVn+BCpfSXGM5rHMle1vDUSjtT71XGg
Yo5zZT4Yy1atRN5hkhk4v6ZZDfCmBNRbsPaGDEoPETT0fMT47H1HTsHmIzBZnKp4+w1zXuFnwjtV
xBsfG9e/CO5C8hfhTlLb57NGeEkEwL7jxh0i5Vdlj5a9ierkmAUZfUHwbOsMbY1pZe2DyasxvyUa
pMZJjP+2vW8fo6Q4GCJxFpD+7JKfalcUNeV58wa1hyQ5gEBDZoF2g9CASY8pdHUY0WnojS7Lxzxe
HbWsqCHsR/TPLapKWVo5e7w+JpC1+SBZtPmLxxp2FjfsdfMU1UaBFIJH+dgLaE8QYa+vb0q6kAfp
tBbVdT439eDF80BXzBhILJbTYrAzaTpjoYCdMa9qB41DT+EswiPvmMvllfsYjOWgUkdT9N88cn+3
EAQrMiGq0PlAKc29JAzD5DSIASkKSGf4VmbLIRkF4aESDX+bLQdTeUi1Fm7a56qnw/iGS+yU/JAs
3pBMfmxTJNuMPmhovWQE3HGokSff9r0sitLJYNu6kVlJkSbVZLgVhOkJhN4O6EwIejKjlrH/25ZY
cWeDIEGNQILDBK5CahyO8bFkL4v+tzfq6V8XFH5Hn8T/hPyzdnMmOiQPhj9lzxnrOpa1j/qw5s7w
QPgtvVBCfUvfSwRoDcZUXAQY8kN7jVTAzdtgfduNo1Au4Tt3Aesp2aj+mP0e1MixINA9qpHxCMls
NB8UVCBXsV54NvGG6IuMW3bW6Cb46CiGvKZ0PXE556cF0zu6ylv/FO4E4YkpQQs78miDgg6oxnF/
nOxlTm2SmamTC+bY4UoYnd6t5dESLjSM6Zyam3eWjVulDHUVe7MVQBVJXW4RaAPiWKSrK8ZD52Du
KtPIk6iVfMKsqBVOl5FBMQbQ4X1ffHJJYzoXZll2xYUYhULFPWVEuORbtP8ttyIFMza1XhevlVQX
fPg/eRoOd63Fbp74hgSRB8BLo2fDenVaGEtMI2ySl/oPKtiWCB54dmZZ4lALrqDKxT7HDb7zQayN
w5VCMy7ksPdrwNFx363brQk+XzlZzfSlBwiA1BGQR2Sm4wBaeG7HY8Wl1QktAlqsRDMvks5taBh7
mPvoFU/vj9yqRSg1pHfXdlI3VKJj/Ny3jVyF9iqTMbluGyowEd0ybUwHuW8TdZtnAM+Bpx3jJIQQ
as0Q9yOQHQIjNjfd8QsMs0L42wHTOGA5FWlPrTpSF57yzLWEB6bEezhFyAQNylhD9yCwXRKX44T0
5Ieg3kGp8yQwOZNPdbbL7hfNTYIBCvJB8mAX6MntZ3+oQ0iVEmI+gaX3qXD/1cIoqGIfgyhX/FO8
C3crn3YPlP20uyG4HtdpPxhPMLksUSkZVWl17dL9epyax4mlnvP1bRG3NilF8WvqsSgNJdhJ0KQy
udIwx7rRVqY5R2SrvyWKk9bEILXmXs2CzIpMTlUp/rgju0Ixp/l27DZXJiLFCHCWPgtIhKx6Vyih
Sfnrb6/+xJ2utFFBYNmqJMpIymNY9Vv3vfN7wgnfZKUR/t6aX9KanVbGocd9bo/mn9wUGn0PA8C8
58WbegSB6L0nypsXvu7afdPfIDbRnmEsjftqP8/Q9lit9aSRu6tdizpg0UWJF+wlQ45sPa+dFzM+
EnexJyD2qQ7vf6nSvxuX0pz4Gr2G8Cv/8AKDzaI+NYcWHsIP5Ln74/+CO7f0G/DkyXqYEeuPVoXR
4ZHLsiUbtEWPl9Uw5FWVQwFcZt613uODXqp/icvSGYrTP9OR7cHyk0IHlg1OD5ojP9Pfykf0kKN1
EcmqiNGfehofqx3rWuRHFYCqjbhXlJj0LYqzLqCpxxxn1GbENlFSUMK6AZGJpB0SR7X+akTs8hHy
gMRxHpeePX2+q0C7SPUE/nWbrqOo39ghK60oJgWZwKVodTcQYCAJQ8nz9pKcVp4pP8n28TpxcLxJ
muDn15e93qNAbIRgSPlfKeI282zUgfc7ztB3lolmlPT4laO+0gwIFmNN8q1FCoJEZiotnXqalOeN
b5Q3Te9zK6he7Q26tJ1jYQAuj9RzKsNbVgKpqQ2X09PxJhf9UgYQ5+mtMXipgIsKcz/H045RVAjj
lADQroOphCEyQrOC3q1JeiyUtv8rI6YYwK8Vuwr6Kp/QhwPSaIDTtwrW89y5s3OEBWCCSzDOGnVm
eZBDHwaX7DO8EI0xQsCSXq9K/XsLjHqGmpR285sAZ8G/wC0vFf6jOVhfHXWtBM7NOBnMCAm1u5M7
bTbwcWxvk91L2JL9BCypcm2BJe7mANHIBB4KIwxSkXqH/GgesKQwJipXa25yUOFM3HIT+YIXCpLM
pKChdi+Um6ifsNLFSisZVZ4XQCnVK+MCrxMhdEd4WlOEiQdAVuCpx7Yo/6e6cJ07g84jXMPVJlaq
Hds31j12nQmz+YHLGUfV7KYenKAaQE8TirsgoyEcaGi1Gubffpi2hTJxqvHWwlqCUl3wZfhzdYNO
gns5U3ziApwHIRmAtiV8lUxCz160ABqDj8/+p0ARBIskzVDPwAIrVptI/NYDD82vYO4nCSTNeHQj
5VJAoOEcIgJce9yC3G+IV+m5T9oFEpEIemt/H1a28pqI5la3aS+amENKX+ro/0OdodFV1+eDbbK2
HdxT5R6QeIjrZeL7d8Gw9mZBZy1LR641MMKotHK/GbeqXGH2DS1zM/aspkjPFtjoAe/e/d1gna4m
2kC3rquRE6FXP8LllxiOZe9PLepqVSj7IlLlngC8IHvoLDwcA/Vio0rxp+5WhpGfyfLWDtyfWpC7
xlVeEqXK6gZJ01gucEZ2i6gpjXE5eHB0L8lcpcQztCpwn4PBu0CCWgBCIezJBDk/434j4oTzb4U/
YRwIiiH76TvMUmfpbq7LsYjdPp3Vhk88X7Jeu7fdbVoUanWqy+2NZlJx50tcL2wil7dYD6yw/NCB
bRXDFo1b9NectJtKmr570ATyLXLyVnGErM+1LyNnBMw84Y9HXF+6TDSRWJQMBuDBDVzpCJ15Qbu1
abqyKgoLIhg3ROXW8G1hTFPM2MKnuEh144rU4+ygdyWAHSfG9dZcdR36HkerOTwsj5CPhwByqh+1
6tjHCF3rQMO30r8p7189B4qaRbsmeUNqomTywJzYI70I2opoHIZSDYH2QF0E+4wHzPQ3hiF42IWN
MwbSwccjrotmmzyZWESzhQie2WkNYx7oQ/j89zGjxdTAAAKvQ+i+T4A9/rbKQG9PgT1FqoR/IUzJ
4Bn5f/1TJsgWGYaMqLjThj0Lbb9XzbMjf+svjcBJJYasMPdMTA69u8d1piwo+SWFT8BDVnuVm50R
f9uuobSE2gVkdtJKpWPe7Uzsk+0jAN4UhhscepS3ejIXb3SVqsBsdsC+LjXsRCnuvebNduu51KYf
Jcn0Bx+Uc8wr8q1X30qFFFdjtaeB6RaKV5uZCh4HddPc6NIb42Sd5T1uUeS2wOCWuzAaL23REyrq
FKVJEX0U4QWs8aIknncV2BkHUQJB3vn7nkcaZDctdTCWULTGIQraOal+NXcJ87XC7GA0qy86CnmJ
3kR517Vmo1IsQHESt4AwVAZb5xMNUH86+2aYzF7f5g1j0vzyXMpRvW20CsWcO57QuK1btA4HX8eQ
GDrJ+ZyywuMrj0Fesb8Ju/f7mnXFMKLiVMI2Ujyi1aJKnXBmVQpaIwUMrNknGJrGUHESNGeCcAba
VSPqTqhO57pDYOr6hzZ8cRZgUWWUOPZLLRyYDJH5n6URivTMWsy2cUGhp+V8m/2bzza1sl2UbgBq
xpLFjBcIgqOcVjgY3XVh1T7tcrVWGeueWyoAUIMXYOicLfcvEKrLXxK/3BqzBWKakHpScynb3s5L
wPTmhPv8qsP7WnWtBxoH2Anm4Fl5QQMZiu6qgDkqVB1YijhyrJ187Ya9FRYf5BPqZ/FeF1A02SPl
z02blwOh0tmNyaz5i1haKKK74Q0fwT5sSIq22YnSPhvi4NaWGnBoYMfPBngpF5RGm0HUU6cmVSLF
ekB1P7z0rIZWS9s69ff+TJ61raOZ3TaA0WMR4n62pXr3EWrwuaB0Uv35xClfLB6bPxSghO6a7mri
nCetKbPiDObzRp7DAaZz5BbcPxvZRed3XpVu2o/usSj6FWmVFtgAmlw7/rhUNCyUWLXND8pHtZT7
F6zpbhTw85vK89qb65upHoMJsG7SP4sNpaD1f9D1/slsQZ8GMyZnfPaFu21KwYPrfIPO+jrjGS8H
WnKuIMlnQZ1GsAf8PCR3EJgKfDdY1z1wNeOpd0iNAuz9BRnarsN9ITU0Tg78GtW0qCHvdpBzhFco
t9W0nwXhagTpMKe7FmHlKvfHGaiz24QOPTCSusTIfFAm63hrVtEK5cMKYwjhxf3g5PvORqEiN2Hj
veb18Yf8MZYv9CR8jL694DpHeX9U+IrQEBmS86Pe7NOwKrMaMTeYz8lsXVbb7uiel7LhT0OK1TKO
TUvSVx9tq2g5Lc4wcdTvjyIBy6LpjKoCRwO2N7B51LOY8F0z42C/gZPZk+b86V26WwSTWnNqt6sz
l9CEkRbTLbb8JI6bR6jOeGkVnSePvTuZ22SFcSyB1JpAfyMnTU7KCOAmTrnzwMkGq8RHpOKz88uW
gB6N4kSifUxXSoZy2SI4ysUrEl6KPsknxHu7Nwh3CqQlfk9UC6t+cMogM4jBFLsO613MM4ZRXQ3o
d4gxtpAOd3tkKMZmZyVNX2/CE/LaLmVuvpSY43Y2bFBBSygoGAO7k7i19mhOCBZXw8pUk/WF7B2k
CsXdXozh0neHRN5HusvVVOHMxWzxqTyg0P8QHSp3VJC7aH+4U/pbIHtJJJ3JN5HE+PSv9mE5U01o
OdN7WfWJ5tITAhGCItANHR6LQ2Bmk8cByf87SWTrPp91idBcrNsQJrevh+2AAUUR8vhhbNLhaMnr
MNHguHlnyJkBBPl0PKtQKm4Wrxk/TIbDasbVTpSGlCgwbpwIrde31FBGX7Ode2ToLDKxjMbVMNg4
VVougdltyvJcCVCTfhrSrZJKoJ86a/QMZkuLtZTmuyKYZPKJkqSfUpqEFVMXC9OOZPsx165CygmR
YyEfYGztm+h4BSSy41ZY78KpcaGXL75kse9yqdI0bLdn7NLqmEd+ogmGqMSRkbx9Ymq+5rQus6g9
HQNhp0R6ER32CcPBVVjUP+PZGU0zW54FuLpWPH3muv6iATzvGmr6RK8sPRu/wV0G0c5/PvjAoAUe
xDRZVj8u2U4eJIFissMh8mmFSs242tRakCjUGdXosibbtELq8KDsd9jXMZCMC5j4ZsZz2PufnOIL
DKwZB84+eAtgfh4TBuOl5blHsiZIfVtI/8zSwDIowleIBiF1a4Q/RVHz+0ceKZIQw8WfrDaDmsFO
vTj8ijAiT/UqGxd8Na3rqi4UI5PS0tMb2uuCDaafFbH5VdxI5QudmT0/ehZJjT/3MLDXqIBLrp/s
9/C367Lf8v25cGcK5IjXLBHpJcouHOl926Ja8UisC8WW+zu4KDDATvY2wqzJTvvD2cMF/ec8KkTC
YPX0s85RVDBSAorYuJfjNMFzqC8JYRLmKoaq7ml5KkLTRidMHbJWMIhE/lbceSLPk46lLQGUak0+
GzGHpzcWuFVvGcXGKFK7lkpqDXgmZwXVf86WSMdyt6pa5r1iQr5dG04xqrQiSLAXWJdoJDGu/yU0
uhsHdG2RBBes6lFQ0RiC2dui94OKdwCEjbGdizWS5EqaFgd00bBFDzQzuIrxEeCndRGV6idZCH/7
q+wtqbRYxAYcRT43xajP8Rb6peb7wF5vMYFwfcuCoiAsmSDJHdLslZAP0HVoMSI5OJYrWY9goA1x
gyuCZ0WNqEpim2QUcxUINwLgpODt+NXFHq8VZ4ki9ulTG9PvbIdXeLl+ny7eQMFYe/u6f/dPuvIc
/3wWUV0bPdRL2/sQQj+hBRZS/KKcuNBCb8Rn3au7n5fiZDRcuQ7QkB1vJYJh3QiySgNLrU2y69DB
8YoeFXcd85jsjyiI9nrHp16el+vonkHZy3UkyZYJwLbfNUApamSwQnWaxTibLbeqm0qQaFl0K5RV
hpj3A5bkhRR0kN01RxLKCw1scSikDw5t60OdIUwtlzIYGETLAJpnXfTSpaUBftJ4eTMrcVH7HVbT
1z5JuhPEJjvaLCZISovb628q2Pm8wqwegGpXPPDXeNoz8z0mTPZmbEoOszWS6gLEB3IXsDdWq46k
qrbd/8PEwIgmmKy7TA/9ol2l+SG2dJBlNDLtYrH8NBzVu+6WVHx35NV7eMNmN2Z4xb+VV7faWESs
cVieqQdxE/YrQ4NlSYl1ZDcGveIB+LhPiMNgQsQO3J6B2ljgOsk+IuilgUr7YeXL3GksSiccyRAu
batqEUPB8p5L8L83V3xTCf4Bx/cvOLzxeZIfXnftIxCJEgkvLAj1+rHZbMGozoXK782ZWaFt8pJI
e3FAmiKSSdhqgX/7C5bAxJYzRA/xSRbUVx25frzNsNKVAYs5+/E5HwkuayX5VrcmJGpko2Ox84rf
3avT2Ij7Ovx1meKi5hWDhjq/LkIcqyVB+xaYkmdOuKIOT8gyoO8JAz+GzNdQqRCMeZZmjwBi+nqg
6h9AkjuZCi2DBF1/yesce7muaRWSf5pA4hZygc1EJuELVud6Cl6LlEy+tN7kt6iKGSKiy2La2lWA
Mu/R2c8kjNhj1dqmMD/mbas/TlYZ3obM1qq8Ifwqa4n0bKIRRNehiDubk7rvrTsKiGMe1S6T1X4R
/jkFov6jBrnhUE4znt8iPwdL2Mi3CnvbS2kCztzK79jusTvnlJDBoypCIRAgYPuqD7zVvpqYExtP
2S9DQBCM6wSefDh2ucD87o1ultAi8M8fGqQCs8JjdsG/MCUlskWLv6b3IikbYjMWilZ/T71f0Rz7
/sWbx2g6OiABnT1/bK9hPVBDa0b4Xi+YMJnwLOfQ/rJeFeQTSSnm04xwew7GuVmOal+xKCYmg/E6
1eu//WNAzDO3+EMgzRuov7dSol4k/j79r7pkCQ544NRGPDLMJzQIlbmduILD7yRCT8YLrv0nWnJ2
bSHa2Lk9te8VG3v33bm4M8p0BW9vbCS6P95un7Jh/kKAa4oY5ory7qURNwYIEyLiHrHhu/EnmGIt
NUxLpJ8FGYk5ImyqAwqOKkSrwca4ZdSeKzkUrLHS+Pnj6D5Srpk2yXKSF9EtHfZt2fSCozJOX3F6
WrpflzHZy1eocB/ntUxMopM0n8/vF2GgwhgGifkknKVbfemOofk4u86q2UK3KjsZirRLvwGmTdwI
cdzDOd5zmZzlVL2I0Lxi0nCchMaPK+EOuTLmZ+Df5SAtHFJcYl3pkaFCRUSD4yWCy3F1SYdbns1p
3CA+xXMM+MeTw/dH5Ogq8MbKxWIJS+l9F7Rj4c1aLAA7TbD3VBWNAxWdWfLYC9uw5F+IHiQCLfpm
bXWV2q8Ru+GC8sf5wZmUwfTFGhPlTqKFZWYAuVwFUt/DcHcYG9bLZYpEy855lyU9CCWDfRmYYz2n
DnST8Utm2X9DRwuYcXu33cFtOy9jgI0mpWrAQLU/i9Vfbxcwi+xBGZ0ukX7n8VhduLnqpPNXzNQi
UszFfi5SEnTZw+3u4ugoQtKoRj+DDu4j4ln9sfu0aWxCfL4mj7sSMLdyGPGhOziDGk8FxOmCoU/8
yZqUOwyirp1XoTgSMEFdgerQAMnu22XLXoH/GKTGdEwy23zoXiD0MNS4q8knawAybGGAJLPES8d6
UQ8bu7ubxvghHfk9FH7BjQuc6I7IWLy7P4ZbrTQhZPfbfOzJJnr3/8k07fvYrFOmTeRhoFJFe6l7
YnCtP9oTmMd8hhZRw5hpP+aNqOwKvM4IUufZsozpMqsq2cbNO1B7xkZH//w8KqCDItEuX3HobJ7y
CmSzeO18M/DANfKkp3dtKRSTQzfLFr35/3W2Lxw0QvIGTtxNEv2PmXyCYRZKmx+0UWCJRYIEIAl6
wx+zJqnghmFOM3j1+Ytw/e9ZF/vhZW4RDDoae+8/odAm6qfUaA3OTtmdyKmDBbkvafvZuiDpQc16
EfW/l5t/MY6OcjQxZ18ciyZmQmTSuNm7+g97PyIeIaOqotCDtc9u/BrCOaRHRwfZxMLt7/0EJlKS
0zuDy2Hl7cP+OwOFq0NeWjMGFmy7PGS0Kelb4AUTsIainNsrm0oSWIRNkEK2UaAF9axXA2Qhb1mT
MoVWLU+xivuGIufNquy047FLaKXA1XiM6RXMKrwK90LIEzWHJ2ryX81ccVBba3s/NMGpQU+L/Ow8
XEt2a1CtuRt5hrQdpl9nquqhukHZi3AYesr8AZhmMmmkwSV4ErKv+2B/Ce9UIpZdvqYaPwegl/zC
V/eGhiCwNbnO2uI/p7OOW5pdezaaRfOOe0ArlSlgHcES0BYA88LNW9TcCklhU6jeMDdv2tIYyE0Z
W/93FQrMhOqxKwUAbJxMdrUXZ1VaOCJOoIxzobtWuGk0dif38f8sz75HE47Ia71J6f9rkxI1EXeG
hTj5HdbHRvqP4PjsV4df0zwZ83Kymx4uvfglNP2rXO9xM7KKh2zNYHLkFogW5ilajELJsJYuubaW
IJXZWbUCIZ2G3t/+j0H6v5RW3kUNfl/QcxETl6u0hAiOaT8CBd9LBPRKEkElY5wPewqn2ZPF+x4F
0YXK4eblmiQ9He/zEydpLSyUFRiXKJoHmLXYUZ28DFPucMskDgoojTho0SO9Z6heAYT7ZzvcZKR0
c+0TnKGw4fxlMIrUiKY3dH90EfNvROH168LVWWAAbb6rpj73Ss28gRKmQCzIUC5z/JjgNKWqc8o7
Eyowq+IOFd7OB/WiwS8X/fF70fTu4KUYsq/q5LVZxCEm85x9FUcg79TeOUppYDNj2p1EzTs2zDUc
Jthrs5skeqU0rM2xuAXrmCo7dtYN/IpOxqZpoXs02cLEKXT5DQq/sTeyOe8Lqp2Jw7kMM3F4odG4
uHwNOhKronM5FDcy7x1GXNMb3u/iV8MLwKmhRDUMf4m5oDvFs0+ys++rAbCOU9mD8u+Rcx2a9yOU
Cvs3ITZV4G5zxZIpLGs/fU9zxuq91zcuCfmqy1lmuY4RoVOT+YOblFeJYVKbW13PwidIGvXlnDF8
CNw3xlGrMJ0UB6ldo5fmumx3URzMMeoF/I544doiO0Ul9tOkf6hpbOo602glpSk07wUe0la64a8W
f1zhKTj+mF5bd7T9Vl4Id002ayQJgfMtPt0hDpbDPZlTgnJBVCkn68GRaa/lHZxkSdCFT5iLD+Jm
pykIAMDp00DMoANs16K4gm6IKM2brNXlNi8m/OjdUy66ailhM90iobsluBazj22VYMXa6TmAdykx
xf+3+pdhfp3uvYUwPNW3oiiwqgPunxrmKCLkllzrVAfyzUXBibbNxoi8FLLPOW0L+mg/LhtUslQD
qmHDahWzgr3wR41GscdsE0tJmDXi55WA3ei8BstpxSa2/xB0Gk35wHGcxHv8R9ziBs14Q+eoU/wl
11lrO4l4mG+nnbhB7rsSGFnHSkK4Z2MsCTU2JKDF5AjRQEcYyS1cvjuknIVbuzlYf/OKozYDI3h3
66If9YXBHzzL7zp0rZprggjvE3OdM8PhzlZjtrx7ZxAwvO5k8ZGMyBadV7S3h1ZGBIYsfYJ8fio4
VpoNk/dmwQuGi3XhsuO8SCRDBFgKcc3DeoES85AhRZ1JjzsCJ9LnGI7h1nt3Zpa5uqgKZRKGJDcv
lIE4BgdAo+cgkEPEFW/1CI8xxlWlckIkzKwXiPVTw8/gyrvdm47A7aTRAgljzDJKqjN9+XLvIy64
tHA9E3gXvyjXm1Sg7NW3NreuVNJtmwL5gegHWNv9fKWkC5+CA38aoE5nyl0rrAaOQGmRarYWfeWs
AmSfVMhzsSVrY0fZ1RJdFbqPt14Ir5HlxcVbxNKCDPVYKf7N+pIWGiYCmm6VgLJ/ovI0lwbVDyWD
gL/RRsirxFKOH3aVjo8zj+vJY5p4wWE3d77JEMlzm+EgbKtlogcDosHqDdmCzRmg1tHfZwZJa5eh
PRTgUs7soLidnB4LP2RHOFkg6OEKFZ8XSl6bQz+kfNF9Jkegq7rICLCBC/hVGznBO5+MO88s03t0
VXwjzQcFwOirvHRXtgAXyAMQfccfPXHkY5GswDdMXeRefavAiFCNrTNtz7SKXlUpnxr/nSF9Iyaa
LyLA94KX4p+Fr5XL+XBvUieKdqCaAvDqdc62X5EvbS4eVpFCHen4+JmWwnZbF5ze2aNFoJUcAzS0
xmm5CztKMAJBQCqAc5GN2ojEXZRzQacZ3fgRSYMNzje5Nzi/fXnvW0VeNvJApri/3Ll7YQTzMw+Z
CE3RGivp6EoOcVFNP4L7qYP2nj3140SK8vX+/Kn+eHswREXMOIH+RYVTbB20BXmy/n4pnEDN1Lt9
+p23EGYwW9JpiS/CP3V2RPpisOXm3psbhdbunfdlVcfc+Fp1DiUUXsz9TCs9e4LFyChE9aaXmtqs
i6wR86h4fHSl9lf+ndDL2OT5TyyVgujzFXgC26bE3C+SeHk9kUPKTsJOilkmBwCkyIQ3bMWmcZa8
tOb5fdeBQYYWFLiAhIyvoZkLnHsMQuq9qz2/RpZ+E2oSYK07Q48g7uGYJZTL6wlF5lXW8qDEQK2c
spFbqMUUpshRnIdCQZLoJW/PiyBfnHrSQp+L9utTv/L6JzBvD7TiEcWfGJWXBUiGkrlRr3xxh4KO
7ivh0WyPmn/Kq4SDgiejuuGD0vvdnuH4SnL+dpwyAYq//RuctOi8xEOtpv0OlhJ6HIrudqlsDhnV
KxlFMlI/SAEtQAm+J0PtUYXnMpB8zv335KwIGmSUTVMKAS7b8Bohw1gHOuSTRnq2qKdICBdEd1En
rocX7dXrMhncNn3eH9oFTe2Plki3PnGQOlREtnzZsO0YWanYOMAabcmnudVxe3aMdOZ7XXz6pC91
PHuGr4VkqzrLxHTyu4AWpS5S5vKuc2WSC8HhKSMsVHbqxQF4QW6lhyp7jUROWgUdkeyzZFP1DfI8
QXdooa5DoBHVaKBmjBXhP/RczwyHIlO++3ZKgXm5jWal24hjM5gclZobi+yh5LgXmDxdpcAX30L3
Qf1418Sfpcp0cO0hTvYTk25u6JjqmRjvHrPRCXY5z2rD9RZTAvoBKKp3x3L7csTGFV4a+AE4nPGO
UK/2elp52jbyFHvFkZ4B52XJREZm0fnK3+glcl7rN0lqRRmzbTF4DnQBJbwG2cfSQr9Vfwqlw0EL
MFLEPCpz00u7Nqk3XRMvTifQ1ruTRpIVYebq+ktVXROuRXgMJPcRYb10mJelIj2AU1ieuJt5/807
GHG56djulBB9VH04CO2FXDDMal9v+D2tZof7WyTMFnMbBflh+x3x5efPPafDvMuTC3m4DW1KZlqL
QeZjryiiFhI3/JkR0VvwRuhmIyeSwddQZA6iUfkDz43eDFM7AV2AYOv+ZYzuKvN2LEAOaQhNZexT
SxO2LE3YEND1ZydCDmj8flbrAMqkrcq2hKdD6f601+XEVbDM9uLOZbpSNRJeEkYB7BoJVtlS1Sz1
h8GS8pkdr2C/MvLDCggNfwYL/WhXNEGlN2Vt8lU83rrERRXgwNuIVkTyXCeeJ7cVbCmNWrKFHAKH
zI3a+cMscvSvvEUDtwS7SDW3gVbFhHrWi5BnB1t3zASXjgDS65yOHpcfGYy2a5YGHBI4Ah9CcTG0
N2UZfe+XJpqHjLD39j65FcVeHh1BUtOuMuZtBk1Vb8JRq/LQRMTFEDNVflq8Tki5MLDPl/2kw8QR
kjn8k5XxMYz9Fm6kVkKVEHIHvvUXGUB7wDg6L/2a1QZ31W83LM3YnqKfSo8EzYQGZNnaVTfsfhd8
fr8FtaFyqvR6yzyANjWh5qNfQleIOKyK2akQMfeWVw1qqsMh98COPotuDRPDuQyP/UTDyba+Ncix
2XH4hTPHVslxOXw0Gp8Plqn37IslKW7WQ3eIEJo58RAoqx5rrFT+C6zDPZ6cbMDfZqS0J+DHahPi
fFY4VtWqXlpbDlQcmolIlpLQG21TbLKgoQwhcjnvjGODeNviIyxQIv/g3ngwrK221XoHY1VlwDjE
wUEFm9ueg2b/pwsMF5KDW7lklDA4pnPzbOmJbcCQV/B3qUobZOC8Z0oJ43VBndScWEL0eeIfYE3V
pi9Tuko/dFNa+9kCZMKQNahykAlq0okhqNL5XSZNkqZv9dn9K5TEeky/v5n1fpffCb/LwxRIxNqp
J3vqzZzcYbNI5MC0uTWkQ7nxl2SSvufB00hdpM3CWcGWWGPm/xg34eqJpKbdgur0qt8v/gOQyrWC
lLPPx6ItQcsL0gjBLL0lj1r9M9sKW2ic7wkyfLphgsOcYe2wWeV0bMArOzb4fexQuT8XOU/wnU0C
PTlTl2Z4tXBMPp2YHgEAqccK0DGvXKLXKOlV29ASoRUK9LIqXPaCn46wKehweDFMqcaOuS6o7876
Ta/yG47/UkSx6Qu6Piw8e/+g2kWNqR24l8aZ8lAL0b2soyORjIIT/r8Q+18DK/yJQ6PJZ+mIhk29
6GicajQcDAe4faa7CaFFuLLL3H1FR8YVa90Boc01qNFJobrB+VtwmUqjNaPkJiOq8+g66EQkdBTR
YNwUnDoiYOwvbr8im+iZdauPEaP2k28ukEHazy6aBW7Ya31oX8wxc6J48tgMH3j71Z66FqjtmDiO
gaEzDzBqZ+tYo79EXXAdU08xuj5JrGWHtJZzPKnVOMrAFwTISM97JQ8dHg8VudJ3N6lgirejAB8z
vsZZJg/rHgG8fIpui3htwtQjzKF7TT+u1kOtcHZi/4DDoEmNynvTHbs4VRttQ8YbS7No5AX0G77K
xxOjtrheGjS3bxfvz6sw7zWHZ/4smeg9250FGjQlMBhn/P3pOj6o8VuDmvN1CiOAf1v6Hl6omxn9
cGIyOnZR9r7W9jWS3ep/wcG1mXHlQZn8QsF0TlCbSSqI3oLBQCLwYaL1xF1Ui3xSYzzGdeLHdHNB
pUGooDUXDoiEBqerEkLSSmIvPvPIvVmZ9qOywi6kLi8HyjdbjNACpqYP9qjKVTsbpwBVMlsggd17
OT0Q1E3TVwv0ihplQtHMS+Wu3TEkZJ/YogJfP2bEvcTWHSE/gJW7zohcox6LL8D6kj6vbPekLmqV
aA/n/QHy+In1acWN5F1hKDQ9K0+JFnUHPv6zdMWskyuQWYsRxlplS/H6qEk6ttdWwpr2aFZ4FwR7
n3PMiU+n3x3csBbBCWmJ1mikq0tYW7Gl6NWXD2Fr9PLhnbjRQu14ASftU0t+8f3rAYZRlUxsEHjN
kW+vPJc9ZWdatVv3ke7nc8UuuiPdFvPgiFZwbTOH52urUgwU7OHyL/D9frEi+eLvsPutLQEhlHdq
C8NQpd/rUnsk53aiBFaXZfMZdYrL0gfL27OcximdsVUWXy/VTMUuxw6fVpo/9ioaMGSy+7OknxkI
4XYRH/Ahx219QJf17vx1pcuSza1d3hsFEjXWS0yG5VAThsmMXsSGkVMd+WegH0m24BbRQWXt5hkZ
KWE+hAEmbTYi1fYbpSjPaAFW0LSBXW9AuF+cLSwyXH6FAeR6J2/BP5MDWpAkRbUAyaIe54Bh+kej
UFwtyg/WpFFq5AZY1kW52vJlCmRyQ+NEbOICfxlZEhZLC/j+olsFiYEg0YB2QM9WiVQ5mXdE2MlD
iyb6RR16i6JynS0Sq/NfyY9BkBSPs1Ov3f/9UTx+FzY3qdMJjxaaKT7xYCqOvDda1WIA9OmQB/kJ
aoYqpOZgF58iQN2zpJH8dm39Fpr8Gh7Crea4SSyA0WUciSJTXMysal1tbzw4CF5nImHItAIofkxq
01mQPS3GxvEu0UapH2BJSEbJtRQHpXFjEyzTFynRvg8/kLRURWgr0IfmP1sj/kBh/slosD6nNFUw
W1GywgjKv4hXeoay+m4AaF7OZUfb+gqON7rOuqevSRnM8h1HvTqwWu5Ffxz6Fw+po02n7kwBUOB+
fyzF66XYQKQWU5LuaSWs0CDoREWkdGWCUQ+YdLeoBStkqho4uygrtWmQBWcBWgdxf0/RYYX0qGIZ
G83USGVzfXZYRcpzQKmkcPEOq4SNwN55c7TBGQUgf9L3fUvIemeQsnxhzMOQNgtIiFXryXeojprh
yEjXeF/nE7QEjprxPX4rRA9XGuzx6ZMRMbr2os0rYl0sQnoEz4rz8LrbmpOhRKQ3gL5COpi/rL9R
+kMDj9wgPYOgcNRoR0BXPnAIBEzb0VkQCi8sVEEHv3DN6VEufiAvaQYKFcgb1AnRZX6BOx8wdF8x
hsrfxgU1AanfY6ihMxb86QmMCK393o1d37vtJkcAp0tRBvT4ccN3/+1bF7V/OBzsPR9FOJRoxhYw
33ORHhGzVAn9DssAT2faFBq0H+pEOVN7n/V4wussM84IeYo+JXAGNJbfuAMODTS26gymsYJqdh5u
/BeCvN13PfxYCYu8K8D3Zs1/CvGQ2QDNT8CFc9Zna/QKSR0nXAPYtSAY1BsN3LlYdbm6avsr1mks
dJKS2SlT9fLs8BVFGmJ58UkJ4gpz8NGECh+X/hY+R+oMIprWlfgjr184wtI+V4DD421L5a4BfSeS
bbTq1IBRGX8l7zXDj4oWQ9axgc1w01iRzMFh3LL3+uSDa1FNmRzDIrSiHeqRSn/3pPDCda1izSoR
jcF0IL7qirpW65hOI4az9l/DcCFivUShTU2cwpjdqHvOY6GKCbQDGtul6nUAwVK75erZDEua9C0e
cYmwnhKS6ts5aip3EIkYt94jpoFeoe/Uax225NjAYYdoeqEbYhY22S//SqDzgAY9KgS0F3KfP5vk
WYZVLU+omhcI9qNR2A0PD48riX2k4XORxXjJLa6hSJjCEx2F9LiwcAhYDSII4hWx59svLEBF44hO
7GzSdoAzwhZ3sliBR7XjrdIflDzZkFbFGcDXdvXL9YQMBDsnia9O2GRfCLPKrR1CdZ1mAxwSWAy5
Es1TuFdL9r+4Qdjn32tpGj08p/15Iafnkh3dWJUjvgkufIDKMj/3JSpnuKScbP+5jyy89Kt3Qjv6
MtFTLwqJ59yzXqE9ZxJC4pRn1g8/7hE6bU7XF9nEQeiB3ekxmc09j6e9wqhDGkfcpNttRi+KZyfA
Mu7EukpgcqS32HcAZbGpETp9JqH72PUcIvIwrlxc5r4cJVpxJQSDzXA2NkC5hMphkSBEEaU5pmNb
FdcuuvssJX+EabbJCSSUGUxkPOgUAQEaXXzoQP4veeuXBJVADpb9HDtV80k/60aKpaI2VqCmnR6A
abmMZ4AJp7hY27u1PzRzuhcTNsTTzR4TeEOTPBOaYs7j02Aqh7UB4gJp4U/PyG7szF3XroJRukAL
NJHl/cCGfETbAr56paFXT5+a1Q0Cn3pV5nAgyRlj8fZXKYiZj4XGFX+K9qxeb6cE9QYmM7MMFptX
b0yzHhpmiHUpze7N4PAySbTjt+nIr//FzHbvriRdppPEuCNbvnhU0Rt34wYhaH9GEv7Arytfq1+U
5kqVADkGF2R4Th1iRRrAkA/LTWzAcFRLQ4e3AMRoYQG+sYymvuJl2j0ukhUXMDM+0QDDibdXFpDs
aCfSrZGQfyY7H/Kk7RqM1xihPhgDiszh4F1IdD3nJ5K8hz5NkiMu3UvVaFCbTcRY0UOhjYSOspRh
EUllhnT8C0eagKYqC2TC5b11b4m32VomRJWWlS1XHVySegxHyczt7bdPycncqoLTs9qoQux5Ucxx
WnyLwC0XesorfBEE8grCtWV3i6O2fVhkh7D1JaB7Hlb9W99jRhpZJM3JemPCSyLkXXVd3o1DJnj6
qxY8dLmByKDWjl2TUO3EdeOHiAIrczyyZTfQlZHziWeXXveo6l94ArIQyKFGKR69WOl5BSBn7Yrn
7QQBEpSGYHBZmhd+LOBmQW+zNFr8c7QPJerRB0u801hYyx3V721xGvPRmofIqKpI2TwhmSSLUD+h
HSf1LSlQvzbow3YexdkxugnSS1GQ/A9QJJhCujz8iDCYsfLK3gv/sZUH/cXszxPup0UHC8bh5nVd
A0RCVyaWSINPl6Eof4zTC/SDM002H7p0FgcExN0PijkETD8Z1i8R/f/XsNFhVp/WhhcdmjGxSwb6
LI9kUx5Gj+EU3HRVhOckvKt6qW2brD7Ro0sdaKqsZRaPJwo5NcUSAkX+3yTOoKwNTHyBdd5D5Mwl
JHOf1hGYaomizY3Cp9sFTOBmJTIbyfQwM2/wmKyaRStg6MDlVE/wPYtZawRyrK6I+sU+jLsU4tzK
cx/YZUKQ1/OJQM3F+qfByZSx+bsY06kMnMiMZlsfBS7U9aHSh0npam6tVWUsjHqz8/tTjcrR3drI
jgtCDO1SRKrXzuWLwoNxdkhQG7ClN4Kay9e3SEVgLNo0NiDWf00t72QnYNEhkBM5hSpXOcdTmEH/
UHZX67jGkpMPOqEwajTh4rSjtzdhHPr/kKFc0vx56HE+ExgHKiALWt69P36J5oW/OBQfoBtG4q3g
mlCjfvkHg+6DGjxT6JL803ooVusbYSjJTkhS3ji2RZlHJb+N1w/lu+6urdW04YXmSAuVLVbuCO45
jsM9CiJGRZ3GD2nX0eGtIRkymF+T1LKcqytF1FqJ/VVHpZ/jjzMsFNrFWYe+7NpYZIbMyxQF8Owz
0YsxAMHhNNUs//5w3hfb2sblkF+bxrFNF/eiyvVxuvbAazkuPeOpNeFNUh0ApD0a1U2jZqHX6OAt
eLSe7Xo1Xw9yvo6y/GV6+SbbRZTW/E25jpVKaLTp77NZDSNksONZKrWEIwg+o2bBA2TyHPSa7Qo1
lBYtsKq5ZezC9XkIwxL0RaNCxflWsmpjw8llXx98iyHzRFbOIquQGR3Mi7vwd3n02wrzZXsciwYd
tvAidG49/CxCp9wX09GwQXrFfCoQB/ZMmod2E8YgCl0n8QO7BHp9JGlWcPNMgp+86wP7vvhClQNl
49m2Tb7B8wZ6LnR0Oj0sYdCrKW3+B5uEW8b5//bpkjnx17H/fmJJJXjt3T31cYbjBcf96Ya8pTDn
6ZkOHOffDHtV36oBWYCPffMUNm5fuWogy0lU8L8eNa8OF2l2Zc1+vGFn6BUKNU8dpKgOSNuN2rzA
CHEZh+hTC39oDSGPZMccpbuwdVW68aqkiYPyI0OWNfM6yGGrSJr97EXuxt9Izrxa/pCN9VnkCmV2
RKCk+bdSaI5m7G13EhuLYwayyMSgGu71WDAwgvwba/RjiSH6asHxBiiNoybFRjryfjaa4J5A5fG9
W8XvE3J9UEwnwy5xSXZV/UPaxYR6tDd0DXyZVJ+RTsQuJaTgIgVsz1ToghxN287YeJF8KBdJwmF0
GVy/FU6IpqNxm15lDaX+k8cqq1nMY2z9+AXVMttjSbCfp/NSSgCfOETvZz2JD5PFUrx1azW4GbDx
ZMkTjL8PZ/ycgAEsTKizJeNaLvzuoFY6fHBiXjQ8uomTVDOqpYoi+IUatldVduHWTI14gOoZlbhl
6T8+wMJt65M1s/coq5hVWX3W0z+aQwnE3hOQF1yKPfKo2cJt6wI4KT+rT4iVcJi8T1HKlx1iHicB
p6a/FMQjCHMf52RwcSR6C3HbFALtDgw6r9FdtsGubwsdYIet/R6soODlIXDpHrIk3DYGSUkpnfPq
HX8v+eBWMtsWxqri8qTjrj8K/TC3g/RyHFvusXOt0Wssi5Iz2Gnk/oR5OY1uiPGpX0M4ydlzA/GZ
IvXHIqiOZ2ogl+2zv6fHexLHiDGYWbpfSlUiUyiBfjr6aW1jBWnIq1RsFzg9QA91bql+Co8CAMO2
Dd3NW4ofJR05jDdVOiBRGXR3M43SqU42/Wf96BmY+SNwXe0HpzGe1RBatokMq8iLvK5SHsHyoo1o
x8MPszx+AJf5BaRmrFy+U3mTv1Sa38bJf4yk2twGWFIs6t7JlTd3fNfYDV42R3n4deJZR8LiB66E
h0H0pmLLw2MGtTwZQnPIXHpKbCWllQkSr5N3ewhA/eZHveLI1cplmK/U7LUGXe6CaeYrMj1GrTRt
Wy7ENfaJKONS2GEREFm3nCQkzm4RP5vpMxutc8UtoDSbC2h/YnU9e4dAJScJy2QmBhuRKUh02BcN
yLAmr+nJNZNyydQpAWzXI64UsmAlU1Ovi1RFlQuH8HT8UDSLSoje2g3URKl2QnV/sfOh6xcRy6rQ
OMFJYW3Z433b5lrHzIJmclGpTfbLkvzvNKn4/+MAoNv28SeZ1SXBF1w+d7eI1qlscgcbpv0qLaCK
SoaDrnBtBR6n9i5bymJIahX29sdgkxsyK6OepFXAVhHBc9j+jPgUCygcJEZtPvNgnukXrpGgHRuq
vh2RacVNIU29Up1GxGY+8VlW+RTa7lRC8GrUypnRCn5IXLl8VRRXH9O9vUFiYt1OAvkLTuGDcHzf
JTTDvKwUiwz57h3KBcxoIW5cpvDzSFSshtW3U3lM5gx0cPWucnBWDGGp1X3DmJL9SUeSO8IBY788
LvBAh5qeOPcQXI1Bb5YJDgIzUSpbmmEf8bET5W59sE30eB3rOYNHda3mDY06+No7rynDvg/196Kj
iYFtEMshRZznnZ+4GHOxR1yF0wybiHUsW8S2dx+jEKrlFzytJyJSyEsPdMqE7sefy78kaXdOVQdw
FPdLoLCzTN6BmDL1XDn7CnRx9PDwI28L5g98KeRsoXKEWE2h6omIbDv8yLqxqSNepRViGPEtQU5p
2UR0Mu9FP1colpihactzWSWfM22tPEcxWQUBvbntO9YJV2ndscZNZC1xQK/+RR2+sY/HHOHS1Fox
X+TnwMa/CQo4Fa/LF7MMVU25Czn/P26EcGvZpNWYRTnzxKO7ZcJMUNWxUg1Erp3/ktrmDkc1Ybbs
X1brSKDnyDpooi433b38RE6eBtXW1CrTxzziWnosh9oeAiDV7Goq/GxuJb63tQf/uXre4X/PLbag
eaeFtGkml2pPvhKKquxk0FdZskjn8vFxiCvL1GI2KqtjeD+Rq8xKaJulczbI+W7ZsFe4gVcjei5z
r3a2ipcs3GvKcXatyFfAEp/xeECUzbMGQ+7AppDj9kxQI/8T9QxMeddE/irPjSAYIsOExlfRu/WH
4B0p7qrZOCGlGFfpzD7JomP45qnkpt29bgotaDgJANGCbFgI72OTpMb+fY7d666ZMiOYOG/cGRWB
EjOeSUlWAyyaNS4+/JwYj7nfwhtly26XWM+ql9ioFQdUTW5lgYYtFNFHxrLJCcbzx7Wr29X2sPPo
AcF/P49qNU3eRFxL8pET0ktkpNQLWdhOFKbXdjRnEHAmTy7tGU3oLs3jpT/rHat5uyN51TIjQilo
Y3uQQl8Jil0yDOIdTd4uZVVq3ViJ+P7ji9y0W2iFdG5B/H9dS6f4VOpfaE5qKsZhQOFqxbpdeb+7
F8ehpA73rKXYidS92cMIATwadz351LXfLA05xoemI/C9W72O6V7QlzE7h0cDGSascuzR4HpH7dEA
+ap7R2TGRbR3yCnLk/M8xQt0TMjQJu3nyoNE7MIpHldxW3k5Z3qsvnrQV/pXsdpAzcPj13WYsOXl
E6iVCXnrtnvjmewnkQHJAF4lRWanvn2tXQiDBApAcaMlX8RMH/pIfDtxhrGoZlk0X/tgQ0GeQiAU
ZnKTlv/OUhRsjUpGtEYseuuO4gO4Ycs2rxmrQsqYY0Kg5wwEQewUWp+giLhkYfmiXifCUfkA3G7P
nrz/M9Q4j2m5l3v7KLpHk5gnSKnTQ5TzYhxyY5kXsQpt0TRQf5fwCqAwd5Q27aZv/r79I4wBcNnA
9o9xllMWi10jXHiI2HBFZ0RnBGfJSUO8gj+cy/rNDJ62bvBdlMNtExC4rU8lxVmsCDuPtx/Tcryl
c3KyPbzI2ZTiPhYiAnVOPnc8MX41J9qkiUd5W7pMIZQQ6StJx0nVSjW4YKvZCoIaKBwhUrtxUcZ2
88PYxfTShSDUu9C40eVDFScgoNDl8P3FpZD3RQ3PtDDpS1pIC0v2KYfhDIITIr+x/3i/FyMFaDIf
+XbgJcdrdXdp6kl0c45U5j5pRDxDi+ZgCu3baQbsmdLnLruhDC6azNUdMbilt7kCZ7EHVemreJiA
wSar2kHYHz0pLbGW5tvtt325mItEE3Mw79CTn3wMSVp/zovEUMZOFY1u8cj2g+WjNKZ2Z82Avr6E
5O+nUyPVpPJ6wNplsKVV3zGYFLnDawR4F1Uuf26z2zDbp47Sy/GxWUmViElYLSHYZZegczqm8WXg
q+Lyav0d5JQsB/bOPLPjT4ufTmjgQahuPQ6R1LFIBuENdqVvjVSxrjAodKxLgyN6ajwaj1xJw8Pu
aqu26yLPVh0HMdEde6tjUqIKdPyEQWo0wthn2uScjxGvyi1LRoFyj61f2pHm7vmQdbOMvP9G6w/v
EsnIDm4NHR+ObvLBF1BbSKoE1GLezXBQnp0tiLRXsqXt/2eJFksRLn6PWAwI2C1RTkdvfUl/RsdX
3Vt4bT5RJHBOwkA17Lay8CU7tlUtPTMDubV6GIRU+XUjFne4YQNhCnwg0IbqY+qM9gXexI6Jce9c
OJ2grG77VJPYj/dgVFw4zH2Gtuis6qv0r0HnTK2kl3vGBYpCLeZzK3yI4ZfsTgI78n9h7Ri1XFiH
RybZO3aA7zDrzGATXu02zuX/Lgop6v0oFsGPtWCYgNIC/CupnvXxoKBYjnL2bfmqzvsxq9hEjIqk
6S8dVHtPBRD9QkUmic1gk+KRJWeuHCCOWDmpkkA9mjoZegHhFQ7Qj6oIxnvn0qfUUhFTQDr4rd07
0AD+NiDqYNMz1awRBV7zJNAzzxmvu+P/rYVXHE89qD1Vmo9TE2ARSOvj+rdI/oPZFNcCkzggmL6L
AbTUmS889OaXQBoHtVkLai0g0UKlZrMMJe/SF+BInA0uMLJdEytF4+EbaGo4wqxoanb/jP/KdEq6
3U2gjDiRG+rEDiNh0rBokJDFZO6Bzn0Qvit/SZ67ff9DSNml/7oZne7y3xqA+0KCGr+5owcDRuO9
834LsUdtixSxwu7jmisp3x5HPaUs7TwBJeEPIH807ome/AnLDvBGCdTPsTuzIKe5jkLP9PgJdocC
9Q/Ugfc0vmWOHvTlI6HaZKNHXYHxWWe1KOTzhCP6HRUIPmvfivVC0E4vr8+0knb5w8AZE0btXXzN
XnEwJUJNY+rpQP9svMHtSQ79u4G1vE2OoE7Fu88cjdVexbxYBWzv7vmvotWm7bhhYqJeFwIuqBEw
86MeX4CQdFRmUMHjNjH5jI1qSMUTpBlEjzFQg/Ev7Tbqz1AomKvRVKacz6I1HKFmH5Lp4ifpTX+s
AyAVdMIMnN2CG7jj6VbTEEEBj4S03VlGafmZVjcgtTKdokOnGy7elzldR/2xMcaRvh36rXh1JJuD
BQBJbXM+eFqECOodIfMjvzXFGf2gz81dxFGup+2ahWDJOkxA54sKMPnoVprXZ5d7rQRBKYKkGy45
PdnsuLuo9kUnjt1RyBP1B8bvVc1JvsBzZdYJM/bR95+9ZoSVocqidwsJ76aPtt6ZacjjEzrjBRrO
KYFeY4In5tS/aHRLfoOacQ6N4V7n/EFr0mX9oBhgLwtK+hY9oMz59Yasvc6Ky0Edjtu1H5eZrgUs
uLXUU14g3EPEBvLRee390IY6QyoJR3ZK5G9xQ1+FXNuDCEMy0ICaRF6UcUk7weYpPXeO1KOpY5Su
qMcgC9fQEhvf2sQo3363r5Nfvqc4dMdmPRZldhcuHurnca6wlLaBbfo2qp320y0c0f/BMGmsEbk9
pLnnIRnVlgiAgWWo7zei4Q7QZSlVTnljFcuXjsoCTKYabD9c8Tqhg7R+33s0mxB7PhWty1A8X3en
Y4gNv8fZ8qAEBo2xetgWV8vcr4rE1Rjw2PwbjL+ugC4Mn1djz1exzXrjYAoP3Iu0TL76iCom0sm1
Xf6ryDGViHgUStPrb1+8xVMAmJICAt80rPs5MU90eEeUtjpzl2s2PBMq1mb/i3XhejYSCCI8sOCZ
qzRbPf62rzZQzHYJ+2PvZHHybCmDCAGUIowlaG1JV/orsi9JXegaJn5yIYYqsW3u7SLPXj4jNWcr
+oOKjAMvwc92Fkyx2iLjQVZbuD/xzsvCA4YWFeq8fdEsKg/DkNER9B6gVS76Hh3QSc7iZ9IA2irQ
Lf+50lfQg5tOyOi+RNCXAY+B2146WEfRH7buxW7Hws+C2TaCU4IKLNF+683NPUSs7TcZRijAl4Tf
EgCqXeuDBKDwQZieP6qqME8XXt8pLnlntrKI6yqj/hTXb8bDvXk11lN2khoXfEZYEieV1t4vKIE1
NHCokOVw7LHH3vl4i7PcH1icv0FsG79ufTGZtj9wHV7e2x5+WkZlbKbC66bzZ4soIlKGPHal+7AR
pBwwhVn/8KFUa9G+4xiJYIbmEF4UCyEHTngy3nQFtQR/5Mc1dRjGYwjlA64dSHbhrLLJJObwJAhf
wF3JV6OT+Hr9n99vQ0xlqMi8Ta8q9g47+LOFvlor1H4izov7kMcqBnndaU5WB/PYnyZViqsnbl67
rrktOZGKqhVKdShXrvlf6+S4g5YBucJCF47gJdAlKf7v2ITrZ5lPxpuN5tkm31FFz99w/EPfeNmF
sICQCuS/RnSUMunLYhG648gFjYWcRcgE7CGhwSAugjOq7ybwYxtwL690vYCEqJeKDBGJa87F5tn7
clISYfV0fero611IN7k8uO2sBUlPFTRoSRgpe4YgxC2v6eVGntx16wJX9DWopTZ5EcBaKE/wPBkv
qGP/SpN2ogFYon5noxK0lvJAEsraC71BpNz9bQkD7IjYpALH6SsgP10OjoLn87zRyUYt4Typg4J7
CG7O6vAX9HJKBZXWZmupUErE3v4opZV0c7ZTcrMk1a+/sachH4jx2Vx7kDyf0oXQC4F4csh43H8n
wknSdt0VC4gPRzKfTZfxbyJEYi66G5tvLRv3I/BOX8xfYUqkz2sQjgmWbmCtvSgevibd4hmWJs42
k9hPxogZUh5uBZAIst9LVMc14mBAAHWbS/+wwbjQbdeb2dLsz8bCMVkNEmADYFd3W9EKaZHlnoVL
wiD+jMRSalH2ZKqgdhSyASJ/yvtFJHYmcEQ/wht/IjOSHE8I7S+CRiWkt/POqh953WeaHqDz+Dc/
g+YOZK0360d5/scNmQSnhFQuhVW0IvjmUiQ0Iq6Qh41sw5aKZGY+EBYA3Bo2JgGBLTtoxyzUrl3K
t2x9hNdvu2s3vWDfORSBelby7nsNpgg/hgwAlNauADal4gvIFhTF/5yETFPUuaqpBPW8PvEZQCHK
SWbR8SONg0DmafRKjHqedPoO6bg1pJhnCwOQzErweGXKeeD5zpV/rwVZn7OAd/GwPjxKkCKO9Z+3
EpgbyqQdK4ds8xlQxhfmBgD+6rDZk0tOlNiyTBCs4OscJItGY00wOR3+hIFbT2IzGTsHMMXh4zwx
8eCDloNsYuKv/pTgD3JvmvsfYPVra6qGg3TDJF/a76+6jyYQVzaZ417rPN2R5Z3ZTJIpB1C0itAz
MaXbAbWkLZHuoGtSkhJ3jBDnBlMelQwc5kl4NVpti3hvCdIDycjsVERNg7TI69la2dqmy1yNODDb
SsZiIxKXGhYul1/5yNpxPvxv3r7Df69PkarWN8Acs+Rm8JSWNqiaIR76V/kMTBMRa3C/YwytbZ/2
0QJlZ31FyWpgGUWrB38/SgLFBEzHoeS0Hv7yTj+JQxNJSPfhzsHmttVd4S4nIZWV3fuHV4kKXHX5
zFcj9qrXvEE/9jgeK2UgTXAdy0M5HdG2dbTGkJInDK6DrDGl2EB78yqB1/ef5GFQjY9emSXtbY0d
Qbhm0hDL8xaoff4WxqyGteJT42fCFxzo3s86gUU8QsmuWopYRkJGq2N1FTd5z6H62up0Iibgye2q
ciABNfJcWD9WwTIWO3ae5qrfUGt2Rg4otoEyCikNGZuBOv7FArDlVXaaxX1hg2oyn/d1NtObQsNB
yaUbzKOyLAt1hEcixqXecm3INnX2qAIY94IwGlyOhLBAa8ywoF15JvDxJ5IRdd1Ns6cfcw4XMs0m
ZPj3+N+4aJZWevqxfK7UP3hWHukyMSTBNQmLfaEPAQCJmFJJILdzfc6HwA1XZ6w7xiC8uE8xui2z
Qcu4lJHCvfzMIVgZwslN3HJN+0jo8IovniODdyq9BJTT2cegqYC429XfcfuKU5HsOCUAk0ESZu6h
g5yLomTE49IKxq/azMrZcKaYd6xT7D9lJ3D+eG6+nK43zuzus8RWENvhAFSVcHW3GzTk+ygmxrsj
kGF7qqDYq/mjO5T7YDl23ZXzojd0MtWNZgFHz4O14WBRyz8MkCn1yOdq787gFDUp4tbuFz2uKWRM
Dc4hdTmQ+Q2L1xS2DoKZq/G7S0VBwft8/Hv1h+9hdyGxrWKIoY1QwXQsWsHt6F83vyuwHWE3A4t6
kYPx5HH9rCHOFW80UpPDF7CxxtdKWYoHDffd4Sogx4/TOYmXZLk6j0XCO75z3OsRuHXqJgQqd94r
2uelL0S8uniA+yMVErIlEei5Lf4g+f1qkD1EvcVHDvE8fgHtv+KS1AXxRZXrnVOos3v+y7tuYLO9
9b+uRZwZdVh6PV7O7L3a8JTKfTqfSKTBS8UncMLB//SGMhHo3c2dYPZfbbf4opUcb9+ACFWKWyBe
9/sIN6UO9uwelYMdZbWAJkZIehkhcmY2ewEMfZG73ihkHU11ESMO0ItKDRH1OBj+RyitK3bA8SBN
1KshiufrRbIiMS0iKTpU2IAAfBMFSJO8Mcf47z1I6yYAYl+9h7pMc/QY1xgxhwQx2r9k857cixp0
wzjdd14w1Ux81NnKgemZ8FoWzsvW0JqrXoEH1gk99Zb3eU26HW3X/CU3BJDuSNduYRUK6ZjYCpzK
cVzl9/Di515SfQheQiS2SJRADD5a085mbL/pZ3zUXEIKo71VRvsHvfKCdXQAcN99PMGXt/bc+kSk
O3wSZn52nmjyKXM7XLqA8aHDA0sUJHfj511b9dMGlgsbzlN34AaB7C6HNYnMAUn+WIW3NL+sb2vv
YKXwpf2U6DTXoedzKsrMJnmmHqdTHivJSdbiSNCdlpBZz8TkBO9X2XcLIJlyUqYI9opNdydPe58b
YVss/GZn8/YSnuf02WZGtfYvQG4FB19rULBSfipTPb1vRt6hrupZ4xQJRkbGcAS7FgMYep36Dom6
wvUtBjMcgaQ+XQ0mI0EwJXr4JXvpJj9dqGMvCICG6180k0kyVocH5rA0tBSpJ24TlPiMvFWMBIru
qQorRjm9f3MVEGJ3lQbFdM7NNz/wbH5SB/J+vHhtkF2QEf8o991jneNUKLJALRPvULNw/1Fd3JU7
9ATLEi8KHm8X0fQwfAGaPawpborpjlz+w95307XmDlygd9w4RpYBOTVpUoWw6UoAgljmRgMysg9I
WycKDIG6vj1akYt19Oxl8WkNufnkYNYVzeg7bnekCZhpNSW+3EHduz0NA9sMqcY/21sgBkSq43eH
HuDD4DVLxQHlJZdk6rWJhTeD6Q0SjhLNWiGmhsFdANqSri8ivPRKEy1++pAPhvFTFZRuXzfw/A3u
rACTJ6IkTVKbx60aaTuHrjirzc4s3d+wrLb8RsiSjstTDe5wFVVYa5f+OBTfVJ4sf76Ar4dTKk9r
2i64Xe1bbrruqUGEW3129syDRex7UPVs3f+e4PPVsavyaPZH1NRuTZWEJejXCybj6AdAIKimZnkw
M5jP44b/EFnvrML+7veWSBzbdr8cGPDy3GK/Bb5k7ltN90ZzSqlGDg6e0OsTzK9KLAGP6ojU9JNe
YFXf7tdRwHc6h+p/JAZkGYgnCAP5YhNNQkLbvUXarjUdF7x7UwUEepooS0SUNS5gyFZcL1FtVgIb
8lE/JxGXBqGHwAlbZszEqeK0MD3WcczXFrxubyzEagQN7CSWKv4Kuingx3Awc3xBW+lkWDchTjnt
oQWaW8gpF+krQilHRJM8KS7uLb2a/66CccM5XaVja9VFRGq/K+T1kvp+ydfu/cVEV6Q68XnlvLzz
AAkDKTmbpCch5j1vgQ+1uHjUBQMxNf5adzRUZCphtmKNqnmvdVqlTiGxGC1f5bJISRX9c4NqTLwj
tDEBLehksqE2uWkwTsLzYFSrFbBVhFlnSK8l58/zax9GOBcuKE0ehhbnkYLBDcX3TSJjg7rsn9DX
Vid7nk3GUu0JN+hlYtZMOWAK/IPHbeDXnAOvXswcBA3Vd99FV8l48vjzIZdWq1+UMewtRhE97MiQ
6ZdqGuM5459H98K39LFKQre4GN3KUZPz+aFNhfy3P9nY9gnfX3ELWfoZS1Y82CEalxeZoqXt6kSy
QtAUaEWG0ExURMYahCPRRx6Un8S4uu4tGGlHHNJqn9nZ8rPD+tQ1lKE5AakC2Xn+Zp85p8iiAmJp
amkrLrR3NPEMziM4l5Vp2LgY207Go+qyIiVfIUNZnOsfL1RANGWbSzNdajX/XtcCJgR7MeBo2CoU
hzj475x0FHGO2S985WEoNS8gCkaxIJq19LQppSK7p4M49pFKknCILkF7gA43k6HUXep2S3stxIk0
C7TVxmvEgs91zOStAGKBobkHiSdQ1Gh/JqcFKgan8QZ/jrZn7hqdkzD5TQmJf35QmRW9KVX9NgB/
VjIr5mVys4KjokVH4am+olHIcWvUUuukNrW3MvLUlyceA2Hrb19SD+z8I3IQvezmqB9LQaRAn9h1
hYLKV2uz77P0aAupkd6szPKVXr2Tw2vhNqWcE/eOsnAp0MkoFmnANl8VIxCMKOUeBgknfKn+kHfN
bMP9Q9yJL3pKxAU+BvUl3udPp47iKIIfSi/ZwRz7ednC4NOYkX8lZQ/8X7c7CwyEL7JAsZ0/pMtC
mYylsGr5jEIRgL2xEQIacYs/evTEvtrXP4xgbAoe+QOI6ANdI4zqKav/xyoImRsJZU1bYfpquj7B
r77z9hVqoI/VBz+RAd8KUU8ZyRnqDGiDDTOX8wFPwyphf1WxhXdzOcFmhsfMwYvLgv93Og9L58ka
A9DTJuJZYyJlMg+DBjIX/HsiJbB7VrGICDNqxRrGx+STIJtyIe+ijYJRmAdVsr0CHqx1x1LIwHUG
CBVCDpFKTQIh3NBHDWXJ4Hmkq7Es2Na/HGrFWDVXV5DiFq+jSViiCpGwicWONoFM8ToJvgp1SjTr
CDG6V51GKlvA/kfRW1/L8zDlxMjdlClAQhRAi2tuaaHQCzBGry5sb4U8K7We5hVgTERH+/QOFctm
8mEQm+5J+VAZNRbeSGybknsxK8ShwdSGqEf1BCNlgAf5iL2Y8EU/X/4cbbil8ufpQMOTJJSH+4po
VKXADkEdNzx2H1gnhKyKtlHn85j33S7kgGX/qxXlPzrxviY56Gw6WpFHvzGkcqjbaiVnMNAiRabD
7H3UGiYGZCxmqGlLB7DilyufDhNUtttTZEzb6XKMiBSpykd+vv3kNn2Ce/bQC0SM7qSNa8lWbNkU
Z8vnmCBS4VXkcLAsw5/cZaf3jHAiWoE8tay3Isof5dc0cbtfkRx2XzQAiAWg7dMP0zBjDdd2JUYh
Nrpg1wI9Q9qrmuGzwHM/JEUXTNKSwTtBZ+dApfq2f5zdzFt5dall6XC5mTEKjVyEztKoQwy+//++
q7QGgZT/8Ce9gdhym3cJLXs28WNq5tPj+JqmqCvgBhf95TrPq6o0MxgdfGqt8wU6icDgqLbZb0ej
e+B84JU6h8TdmQiwL7HVbWd5+D9BW7EgzEdwIj2v0q1jKg9kO13kv4dAzEBfXkHAWDn+83AHtoNy
OYZmFrFlzQ9r08NmV2jGOCX5kajnET8nTV3dMG7xTTPSK3YiPp2m1vueeLxh+FPkkC/u9+XQZ/jg
oF8jUUtxH43s66LUyjMo/rfcCd98n8Q5jNVUgbRB9AqLbfjKY8C0lcaEpo2UBViZw8eWmW01iEpO
7disiOHavF7jRIm/zR0rY11lHGcSYDoRhvma2GG/J1p3eTWx1XqAS7GK1vBmghFRdPDdBr/jxcxR
D2n9npHQsMdazPNt8T0L+geNt2L2G/qYuW++SrXHCbNjKkFB/XMmmt/kgzZKCCea6moHLJCrnPOA
0RH96V0IulETeONzWhro7yEkzJt7hcySBJ2kYO6/3722kCVjnk2P3+h4uTA6t5GuiA7oDtwBcG8l
3vLKheWB3z9K3i0VE6UX9uTfxiIdbeu40mJZmAOch1+z+8cobHpbgyfiNK+4Atlgf4cEnVbXk5e/
pQTTn+6BZo9ujqVpE7WaONgs43XCbPn/Xd8YLqDl4uagAVIiFoAWdXR5sRMe/GqLewA+VoUutwgY
fMV9u/BmkGZRabxgH48csJbxe55uBSmKj338Yv+j3GcTMyzS/uY2y+beLneaYTV6C1LNeuV2kQVw
EHlYBSN+KWhZ4L9ZuVTzH6V35C3nPvQBM08yLNlbaIQwXXfm9nOFr8DF68DsdesUbL/eArc/vU0f
J/OmT5fBBbBboR2hTDAE/4a3iHqyqEb6OwL8KnRErb9u3/hp07y/xkJR6LA5Oxkbqm/fMcsLbL8z
5zvVg+l4RCKztRITMkhz+i8TRFVWTlzLcI02yJZOMYwInwZcRJRuT72/mwJtoiO3W7d/MLGsTNw+
Sm+LLjLJfafrVDcvDGxNvlxRmMwWGV7B8JyJuiM5Ef4TyATXahs8x5H55y21bJDJNio4tGhoZvKo
slPhO17YnFTuMPcF9IgJpHj4W2ZqADxpjGXy0wCV6iBWVmdx0Cc3azP+xDGYVa8k0ExXiyO3gzjG
NC8cXsLjsXpnjw5h9Rz181qAm+GPvkDHcTAYRF0RRTJcIGQGAHNQS9UXqjLZQ4x0vVgyZlqvrTXT
/Sa2yFrhOmPjoWDpuiIPkOx0nJRjhCQYf7Un4esBNFBT7Rcd/jyjygLp3uepWsxW33DR1M+yRzID
1gcm6F2lqC2zby3omojTa9DSXai09UnvQDDsjQOjN06fZZNRU55gAaeeN+LiC77dPfkP/o5co8rg
wkomMZrCJsfO5jO7mt8A555fZTZAp1hwoGO8bWGH+7hWbLhhDFyREbvsmh3gRgGO4WYHmNqc++3P
cjUb6NUvv7IeIrXeYbuyaZmVUbv1cLJgypdNTxS0d1GRivEL3+yYA/9eP7IOTdaIlnIzYxgU367O
Xii4V9g6mtfbWkFI9H5TTT29INi5FlwTrxH2dsKYdilJSsH+IDBiqmm78IvxsG5u5I3E5eYIA9fx
Vhv8+M5vlm9EMT/Mb2z6InVUzUbcp/j3cIlick5vgdAFlSTeVOMUYaDom7qpI85EX+hyzP4mq7mU
57c0G7bGi+RbfP4rSqsFY9dld2dBf3yoOE2+8EGeELUn4NRQzQzfUVCKuI18MPB246bWdjAjp6ws
NFjIIRKT8ZjHnFg+9NqD4gj2OiakNva9TzQ0JiuJe/wPPM47wtTWkhQf3Y2Fqifxy15/jGL2hLOS
EGWjtMvyuSxcW0tw6nx93ctBRWB976x59LcUxrzeeaZDqx2y6UzJQb1QgFmjy6N2ZMO51HBOulLh
4t+Cm4FNUBMohNVgWQcu8ESph+kGmGX2OmgG5DJqG2Wn3HCQYH5oc0wZ0ZKDDu/F/B8HkAVqmz54
mUDwbC1JbueXeF5KaBUnL7wOZ4rxcD3jzzgn+cLw90nfUQ4XJ35T9ZHT+LeGgkZvzpemBywmIfDL
s44qa8bXK9MKl7jNlYR2vTgdvyycurPiIOtt7Ar0zYbssC0mIyHR0Wn4QYoxJZPldJd3JZHqdZ+s
8T3XNgkKDJLG80+beATZIQoagaWlRewvBfb5VnxiQTkNhKKI5bsGVcJpBZjRsI1al4R4uICHg8QF
I2zAq2WaA2zv8900xGAS7Y3UERuayf2jmBkdco0ZhMG8KT0Ew0OoxiOwbBO1Nvj9Js0w3sLDGSSP
AriQnSra7AXpNQmPdKHgQ1vZUgB9iojsg3q0iPI+6mrA3Df7vtTIvQVwV8RKkDrbtld4mUAhbAZQ
6PyFqaOQ1+Cm5MabmhBSfYTGIPwmIkgjMNzoyLPBxVsIdCwWLlWzcTUGWCVVTzXPZOmafwbL2EfR
nznFkupRvY7pOBA6aia5xHuvOFUAHt2HUQQiIadaMDjuUGBWWaHUdvhibpJ5mjlNh5kMEb+EHhVi
R6TFkGquf3fEgWtQ4xqf8nopILrBHUiQz+KFfhQ+RyEFu5nhTce00OHoXpWNqhpZIdaqf2FSAmjr
n8nxXv8+rRaTpSEN9Bg0p1vqivzzAIOOTcXGaasIJIMAoU2ZRNWTuQHqpSEiJmyZwfWmv3SOGg8F
djSzCX4Ik+6ZLvaNin5YPqNv+iEQa5Ss5iSyEBwCkCQNEj0QxyXkBIPZQU1mDNOlxcGZYJ+cGLJF
HH/SNVRt38o02YZjpgcEi4xvx5xk6G+t/4VQTSHNy3mLmMKTTqkam/oUG/BqOmQH14vOkoSCOdYO
Md4an3LW5ElLJqDwfq1QOlzJzciw4Z4ZGC3TOLtpBA7a2DH6MMIqfcZgar/sNalj0Z7LTpRtvgJt
x4h0lPzS22cDb3VIvmvOQFXghyBdweGXz5Cc+zzkfOQqqkb/ZKJi70izWaM3u/LC5znveRd4tLR5
tmngrQHniSIYHX/C3dHEzHO3vZ4UW/+sU/4VWqoI47wLGMMYzcAgPRSxJ4FroGzdx4/XzCsWfVgJ
y8pZes1+6ocTW4SE55XirotSBnf+YzeRXt2IqFH0imfCRBnixDzquI/052M4NiQ7eXc63CAy0wxm
sjWW48zUCJ0rnGx/X6dQ7PdvkAHidFQCilvydpvAiiRrjakS8T/VlSCAG8AVh2DGnC9Cwa4d7Xdc
WlTUOayR9y06PKD8qK0dMVRtWuzgBsyhMeAu61wT0mBZVCu9DNfhblUwEkZcrIJyx8UjEi/yCrCQ
BVjnb/+oUumtfPpa0MCb9FpT/f3eE21njYa3ev0m3FmtahDKS12KnQVqkL3EXk1GjZ954yPFIAkE
QB6wEVLO2OctBjiT7SBGLlqKrpEa+hgEW6bVyZlRbp5M7BVxAvyNusBRmlXWUl7SdoRDW42TSV27
uRyP/vejZ+Cpn+gD/sYS2SpShDeN63McYnBVx9EJnrqUotaAqvL5UHWLBx4/xyQZQYBqkp1knk94
4pWQxrJl7FwPlWyMusOkrj7mELrGHD1FeSmG0M9vkGwj60TYfsYTz9NerHWhgU8Wx0BJZTvjW7OL
GZd3hgAOcIT1mY1UGBMCAE4FMDK/FPSm3rkGCoI2BAlWfiYLC0/eA711QDD6PaKc1Z1nThwf4ipu
5gc83hbZDnlPeYu1fbQgEJLwgYYAjM0NRVwJ4OiUj9n/+RmE4VCl7Hf+RfU0C7OU7DjxFFz10vYO
HuNJkrdESMfVdNwiqTXxkrR0XYB99YC+7CKPlkDaQD1Xir/AhJff9Lgjct+E4wDH/T6VDIg4ystK
i3Y9NJvAAgAOaRPG5idEcgztNQxF+zd+aStf14XeKyWzL6q4dI9Jvu6v1DckQIzKcBOydopNl/bb
rC4LS7d0R7b+wEJZ9dosiLfQsczUsGbsxdkIQ9911RoE/1DPiX3s1nLCMJvYs1SH3IFzaEjqWpYZ
veKDpo4zoQNXqvya7il0Uomz1GvhfibBABuyNz5L6u8fuTZYWHYI0CAQpjdYiR/mAifzFTfymztv
CYL4aTwBdvZ8HEy+vue6CD7vINvCOH82NMu353c6tjWefRenqH22lUypnVLy+Q6o7P3FckMZLDcI
1r17GdLs89AEbvYpc/EdNq4EtY/W4BhvQbRYEJiam+9HRNKN9Kwb2KNwJHRmejxyrjM3wJ9Rw8WR
0ZFmP8UDM6FWqdaxZF8jywyY3vcmZMk4P1hBtE6KzS7mAmI7IedkTzl8GQBXKygNnBnGSrqnpTTf
ai8AXjg0EUCPWU988sZqkoj7JAgSNSxGyVGwWCHR6OnJAFhw766flPkgUCjyu+kQKaNx3Y10tFJh
7lEB9ZlrQr6GhVai6TbmCNGUHGVfGum+lFh8O7GXdw76breCp7XXeMZpvX7qFeKsx01COu0EFdVs
J9pTtgNPg0prrhcPb3NG+Tf6Y/2RV1n85T/0G7omdwfDOlPGoQFamUuwilW6feeYnIJItrQw4Iw+
JEKTYVBMOJZguIlnc2laKEHsDziReXKyQx17otifBy83pF8+qF0DiZaRpUn/V4xTt3dEaJLDlEJx
oaKm/YQFbuX7dFf6tFXmNq/FB2RTF5OCV4kGoY//9rlhFHPCLUf6Sbd80XWeMpqbkk/yaNOj2DQu
i6WgDT/0mghUAt8a0ts5cW21qE/frWtn7TJT53HNfzMbM2vOFoWgP/NeBf8r/cYSsw/EyjsGX8q2
yM0pWtknOB03vGmkWR65eN2LAwDUr+nWAkA4WzlSu0q/tJXcoMBXYOVy9peHibFBhQ4YvXZ4TTfY
guXNTmwWgOXHvrQBM+CA6R8eWyhgxMFVwgoZJqYTTYBos1yOrMW2nWD1D8zjzySs5aoUOiO3pohg
UCeM+wXom5x/F+yM/Na7okftxqcdIPYTBpneqSqx2eO+YapVDo3s9N9Jr0TrqFlD+PK2Z2lkL1fh
VZ2D1mQC7AtUBwmv0Kifc3m0QVGjUiuJ8d9Lktvd1n0F3CJ2/SZFQHhVob1L1bB/1hOrVqS/Fqnv
/SkFq254NSTQM1uwhoJJwqOzJ7IrpjWE5g41bQrTE0OwTB34HytrcRnCTrEN0nlT/LqdQ0+HkCrJ
eVjd0PQZlyKVPli4jNqIS67SBP4apnsNDRsaYsl88Uv+ZRQKTPwIOvgbGwnhcFsPknGcG3itStUx
ThmqAWwtH8egFBaQQpWgvD0wlNpimXO4ddj7+G6WbfSBwLQ32dIQfW1S9u6pO2k4iruWUAKHNJZR
T7kNCJMLvDRgST8/p6EliKbSubM6AM2PtbAJmkXPYJ+xv/PCr1N9Vfiq+uSorka1SrFguuaAipDM
MFp5w+UMXpSIClvlcChlspTao/HavrSSZ2wlfgqx/T9xZDvb/De3//+S0Wmxtnhp8pbM/mZPG+qT
TkEvKZA9uKEiZO0R5qV2D6fuv4KwPQ6YjXzLjVOOQ625aKKQzxOi3obJTUZKXktOiVp/SVhO3RlN
Gub8zmfuMtLkEhZQhQbRniLgj7yPf/OyAtB0u4/xeG/Eb3iERGyNZ07s2RT8LdSRQTOczFeQisJj
e4iv3vPxex4otGpMeCP3/cgWwfxsOvNPoPK+skqzrWIg/vQUnDTx1/ZTmC796pQ0aVdfMFu8WLrI
r2fVA480ot3U/U8VAFtahrFQzoP70Cp3jhdruyhF2TxT0RJYnV84L1lMaLBReEQQ87su1Uaqw/pA
l7LiuLa6SegmjBr1naD/m7pTEs6V/aXjU3F8+PVpeCxAE/ktfAURt3JH91+9ClERSVwQ+IZxvSce
BRybhBI29VVyAHT05TqTrC3L4gUYMI+If8nXRRCeQk+G/ZmZxMw7LFobaQbjlb7bMS653mxdYk8k
+mkx/2ZO0c1X6u5nE2LCCVZRyWkURos5ase03iyTzKwsUVJYTE+cwJPqFmo+WWXypv416JIoEibE
OL4a7LFfNlzut7g0+uCr/32RGQY21uNz6+0R2Biz5x0o5sT+2xDw94ip6n2AC6kaLUMFUNUeNuq7
QDWPcdxIlG3cwz2XAZUTbJnKYr477UuY6ZqBeXn/WPndrfYOvXbw2r+VhcwtDpeiCBpYouTOJb9k
4TKnMXHnzs0xdOCcrO1V/pHTulfDhfFI2mKvy5ZnU0t68lCeyYT2qkqy1sr0y8A7viEvU5dCIpii
NqwnGip/gMU6yFim0RHryCvRARjMx6ZbeUroxlNUKENHtNeHZF92d73PUFdAU4UBoZMOPdP31IbB
uRtgH3Xz0JjDTFI/wCi34PxHa+ucLGz20d69hcy+x4xMWNLk2WuUltgAKsBRnoJRpObO27U2ikUH
WcxQFvSGRBAlK6nJj2QXI6DYAruLcxgvMoHDDpOu3aUpCsvtQ2o0T4p6u8v+94QeK+yw2EvNqunf
DrrkB/0aaGghCMgZChXZQJO8CilutxR/FEnzZQHO6VQv3B8Td49j9Xt4qVOSxJPrBDlQNLdua+yT
kHn0GX2cQU0fp8m+SWzcdkD1zyYact4L2VDcHBE299BFCUlVwrmuy0GNrokDm+EHQ1378h2qgUY0
TT/AfuZej4w8m6ydxDc8hGgfidvCFciXOxrdblZDBDcJuw/FNkQImFk/6oVTg4mTsP8A/P5RPa3l
HBeeod4XHBjbwbwvOefXsQaSqgSBAuSBya2UmMXU3rKpyli+T2bDSwrFq07T8OrfxF9BqoNdu+te
cA9kyp3cgRjQHD6Gvi24gjsHKjYuf5DotIrdFZgh/086MY2AzebaKW5x8+qA3Bz13n5m/SWE5bEk
X8yBzOoFjmGRXp7IPHP4/WI3yvZvdTSF/MVG3JxhaU+R+vL36utzoa91Bof9mI3+GSQIuotF2BaL
Gh59gjMGgW7rqFRC2hft60QX2nHogexhkXzgYj9Cj3MyOTOAcp+Vp74cjTESbbih8q0UbDjFfUxW
64qLzp3f323Gek+u2NyGcQe6BQNL1ZKhrvJ03PLlyuOHLWQVFR8/Sq6pKO2wPeKyeLEf5p4SVSxc
sniUfduoMMjXjSLAdOInJIHApMufpYRjFCVm4y0odvCV1UEhpq0jc+EjAauRw8ksrE/qVsTFloKH
gBk0WKt0BcPM/zW84wevWk6CaF4NwPQAetXH+3s8c0p0oEOi7h6ACVjcDRB4WXLBBO2Opvz+caG/
W3XbsTTM1G380qmRlQ7e0Pf9RegLmQ6bKoD2zxCaEEaC/6DXg/xeFJLLCqUXYQ2uL+k5UoW4+8bk
OsQD/tCEJwclkrvQlIQ6Swwb93Ac2PJpsjNbgU+dTqnLZDg4EmihAEqmfOZwv9GOZgmQ8O0zYnxY
CYcay0x7unvRmZ47W+fFbKt+F7np5ofzD4mKTGc5X+814vkYhWvZqjp+xXTPjR19L/KKXnpAVzXc
4kLowZsYwJ8Thyhz2NzudxxAMaGkkFqzXpidFJKAv9idOquaIhPfJ6tT5p3RJ9YfHVOocuzeuXW9
5X1juk7ZJQtDT8S+VPqIwVbT5QO4NG8ofihcifNTbsyXDRJuHeIU0EzPb9nTH/LZefKNBaCy5Ofg
D5yUkZPqZ3OnTVZxslpC28SBxFPPFuBzkhbLZ5LvOhpySLd9bk69tlALxVVhN9mqlnxd9lh5GPOO
YN+phEqk8spEXSNC8d7PzX7TDPi6dmJi/rIIzbNQXGPAXmcBU/p2vDa+TeAwHUZ9D1MTyPUSXFax
vWMpPmV5N0X337+IagG1umdlMhjFi+iiNardDJRfphvGVRF9Ia4CEi+y3Y726KOBXB4R3qF7P8bo
hZ94qTGnxnyftMWWfABWYxmpOtv22uB+oiRO40fZliEtJP5dNoaOz3DhON2A5WaIs2IAVmxeMRYz
yqwjhKlpw3/ovrwp36DOqjWfwHQdCAaeu1LwJJdvNbvoA4Sxa0LB9Dbx9OMEr/oV/emgBqfm5lnU
lmvfRp9ZZD9sXCYjyCgag2641s3I9zcGcvxm3Wt4fsO83Jwr7EkeHqWpHvwVUFyAJnXfE24ftHgO
2IEk3Dk5hyulHuPhq7CbXIA0sFZQjs6XQ7Z9c6QX3EV3nzCUI5lDg45CdFsm2x6b28PzheQVfHRw
vQIlWg0EUoaqevYZ6PnEaeIFTfd08OXJa6aSCCbWDZU1fZxaqv/b3XLh1DVPOHJSjRHxlskRcp/u
t0jZx1A4H9pfVVTQE7trlidR8iTJl9HWk3XOLmWpqkxUIcZTL1YWEM4qkqt60nQTo9T52OiZBOgm
NJ0l8hLH27Gnc06TDw0jxNnZdRDg87vkEvpO0HDGsssJyOnNdwgBaD1AiDbR22bFwvudcg1CaDWh
z/SdANJlyx6X1x4O5l888N3NHCjLaNvJsd+XNpFyqwk35oAejoLPsW0HdiP9wwLoHLSdtNji4cB2
iNathjPWuz6pjfzid1gXzzUkC0GC6up8fJ1BkHK0HFUtGVC2tqAzP+GQkjMy8waYy3q3nrmzLDCz
5tbUH3525jhgmr/Cv++3vW4zy32Tl01Iedv8S0v/zaYBgKHlZvF48BgjcQ5jgee5sLpYgdsHpK4K
uZrLubgMUkV7k38fk5CfTOpjHvUV4pfaDcPlppgSRKS6OrTTCwzA4xsBGB8ysOjZaK8FDxUtgwQt
8/VP3kiqZeS+Y0PBuNx5hgm0DhA7rBcONDte7APShE0VG+3Mt1nmRLYjNqYVGgmBFdYNhWQAb1gQ
uqYNWY+k4c7cuULwReN2yP3uLY+z0A74z0zjUyDWdl7HESuX8suFn6hVM6000bxi7AzrOyRWGMNo
CyBS0nGOmXs/mHlsCX7buJwmheyZbSRdIuhrb+5gUYRPUE8EkuWE6hebDEamyPxhhrqlPcK13dOG
7HS1avSDTcM0QT+oMlFjUcP/L3EhtCm96FNUqbykHwzaFeH/7f2Uri9tkkhwOtji/CE2sGtBPUga
37cGbA/N7bEZJKDqHX014U3NN8XFVXhPHDPvlNeu5UYMT20mpYv2FEwcka69TJWAI9m0TsEOenim
JDK/SCG4JAi7xDskGXpxVhG0r4i/579kuq83RmETmFgjwA35feXrWDG3LUwxsJT+ensafenD8qUZ
3Rn5s8VwguPIyAYs92qeqlzS5cwM44tKDC8syvngA4ycebDhioNoEGjaVyyoIwdFyNVAU/NfFApW
c8RlQcC87eR5993F7GNGpMf+iqT+b1dgWs1dWZpaQzNJesaAgdPc6GQTG/c2b4Kb301ZzvogCeOt
qYLMAYobN/aL0EIUoB1DKVuEKPUnUpj56wvUe2KLDv3fHqTG4u37EQ+P61NWhT13pECOxkOmcQb9
o6aRBY1y+rNSFitJeIqjwsgmgS9A/KIW4KGHxDeZFE9jx+NeDtU4HR4O5kPwL3NRcszuyMW+4UxM
6vKsovBFnp13UOykQMU8ZwyTxRubPl63CaifHtkloHqJepVrFhU7ctR60MSg2vo9DyVk54fMX//6
02oj0Q8C/tMFqHlT5FVEb7k0cMi/iMwRwQcDxgvmHPGTuyMCbsPS0DA7d5G35efi+c3ReoLYVAw0
Jor/XCl1eWiRQTlzXuC8mRibQRDHvJKxIBZ2B5KiKzBkTwuyMBtpZhYRtTOeL9NNp0NpT9Sqk42j
7A/2cSyJIIHoVWvOw0wzv+SokMEHYZEgGtu6eVadsOMVrICs8gaftzw1X/Y61SsXmm+QrpxP0bk2
70K6yNOZSOWOdS8/2Etu91m87d7sKfgzRPnN+Cj2jviOUl1KLsC7pa00EfDGY3DR1OihkFd1eHiC
mxCY8SugCmzuDbcP5rFbXBA3oYzg07CcXbtHfNMEONWAvpUWU+kIvohzz057N4+cYwdJyUjyHzIK
A98btcr/aj2XtLsygkYczfkCqJIlqoTmfCnDDdWeNrF5lUmwffTDot0TDGf23iG77tQHQsOzeIvP
x9fugg9SuDSOqIKlpCM/s0RO+1+5VxMmqLxhvQzva6JBefXQ+si1XiJRWeBZx6W62gsIpB8a0ljg
eBK2X9driXyacx30fab2Cv7CrxHSg+gGwPAdC7UHMHq6MYYWFnuu+0aARt6jAuCeF8bOV1AM1plK
t6jqPhFZh70Y18CaKzThWl46SfI89T49F+CNcafq7K/TSkRseQnOoQlnNSis+lECCcUxerRgEjfN
m97M2l3jTOV95QdZvROjqXG61+lvQT6humIXTKy3fPwkCKsJthby5LOagv4SDWY7ILvFH9gbqqVy
YjVFxLB3G0lSuakfIB/mOL/6hHD09cHi1Z74LZuhqahowBrcdkeoV4td5yYD7gPtmJJTpNmknddN
GiH2tXvbBJniJ/WMK8Lolyq0rNeDLSdgFukhxvXGbIvF1sh5ZYhMXxY8i7ok5En9cbGd9wGiQORY
KV8vGpPE+c3/d/wKAE5ifYERSWYK1/tSFLrllsfaeeYyYwG9e2YofpO++Fa+z1f0UxujcAdiAdWz
w4dioWG5oC4lpgUK0+KW58ePmRqn3T2JeaqD21OoYO3bMaK2npy34uHjO6k2d7L/5O5tcEkZ5sDE
5uCDztSLAMPJMuSrlitQ9gY4MS3pqRlkbueYWW4+XCCAM5Z3k8ouoB+wtPw4FxqRDiGltbUD3XhQ
a40iPjtIsdnEL4Ekfj8wXwBZv/qXdsChoH9rj6kZ812z5GwpbvQQEw51kkvL4LwfgyCznvRvMRO/
UbV+QOdhY21MSEvGCPjYlztZyXbStEex57FcoI/W7/701inrBpVZ7ckygKVgMkBpWw5yoH3RflBK
3Vh7l/PYJhqrZcG4nyKvGXgxYpdCV/HwMIBPNFu8yFcwNV4pPDwz8hHNxGYahARBLhkbleADZ88+
FLH15gwwTwQAViFZoGt75Fv8nuKw5cewBK9j8PKM7/srD4tmcxixGHVGAAOkam4aXMNwhQbPArCy
k4IIx/7CXA0sfHXcLelBJ8n2cSKvxEJVzi9SIfjJWgWiv/rfWwkEpfBcmNjgRvg1kzRy0rP7dwai
Jj7dFgnL7MqFQvC7MX648GB6uhEuzjfTwjcFYM/QPdOZKpaMzvAeG1KWfxEFHRjpcgn2pJJuT14O
M+f83ngNHzWEFAJ4IOKQpphop3ZZcWZX0axOR27qrQ9rH3wRg2qEp5LtAv3pdg4+lzvbo0w4JEzS
OGmTLqjyOk+CmxGaXuQY27mBXJRcc2RDapqyMxHcuKuJCOUP318b3JMUO86OIy4toB/lhwQdazJx
cOOOObq6TKnMlFsrYgUjE2VQJ3kpf9b4aBGNmd6SDEwPzsbaUhNwW3SEJBq9bSByHti8F4+xEsPh
cN/RGVgJeT/hrq2TAWR+W80c7nrBvCuJlYt24NsvhOqoC9+YT8BZUiarIVojb27ty0KF8dOm+80s
cqORxKHyr8HriZl6MQPcUOGYbCXAmGJkXpfKFH26N7VGemnKIFRSka13vXs2azJTbqLm2Djfgnfz
EQSGkBJqfE/sadxLC23DdDSF9DhRGS/FiJ+bKxylc91i2a4ElKclAQTfPpoLJHnJ1DiyAFPoB5Pb
xeqGe4a4OAy6cavdlqud0NI6TkJWdHtvUFNaM2RYelheFy3/0JF44gJnvZcSWnRcDVW//fUyKavo
Qzqo0/AfqAiV1XEkkqGMJpnujUJlLWI5PiFrdwE6TxbzO/9tuqsNrA9e4NLCfTkCtcV/jIAeTBw0
X5Q+DwoPxF+6nRXclIGaVz4A/JvLSjFkFPTw5azrHKzKK9zoh8k3hfndJsyExXE6yTxzFNIy9iNv
SXSQVZDMv18+8z79epxIvuukX8Pq0RpwBKJwolAp9AH1wFvt/i2OXjhkO2UhYb2Uat4a5R0gfjhL
ymEskWiWwKgCddvnk3SKy1cVvv7x5gwcFtnai2dZkhP0OyMqjCIlC4NW5DawWHeqtLiwnIMsvmKA
0wFLIr3hUkaS8lmfi4qR5VvN8VAL71gCmrAaB0aTkSNw26G7NDWdPIc45D52ZNHtZVrDIFa+cxBL
0hIzfnJGFM4BftNDnu1w6e1l/zlKH4YproE0CL6T2VsXmPJnpUqyVfydaE/eEQeD7Mr4BtCpbRfC
g6A2CphCtLI0TMQlI0mr5V+LP5msBKBxmpdPuhOXbUDts4eQaNAj2mMk8Qw/9LKq0V290Zt43UFZ
TTsLXmFx6glTsIw+191SqTIiubV9NR+m9aJZPYshIL57SwpVLvsJ21Of9/dEgzg4hSig3I9JgA+F
5j7YP6ujdyJOClycRxdp64YLFn6mlqJLmTv3t7hmUZiVFDmTNzDA9GzbsqCh542kL49P23zHBpmM
b98uqGeQmrN0zNkbeL7VBOy/xEZ4Yy1wTSwRgPQWAeC2TfciruEuajNIEzTfTJ/IiZHLMaUuPnuR
KVqBdqFtlKZjjzkxnDV4KkzkFWnBoJI8htKfV2AcWk2ioBXZOgWEE4ayidcCJ3vAWon23IXRGs3j
GUNClJTFDuOXUKKNaY3FT+WAHoqo4Zs3yDWVm6GMx83rs0OVPiw80CUGqBhBtv8BN9eBPgmWTCl+
KGto2jiiMJxNI7sZ/mk3wmmGWXYu+0E7nf0CCr8kKl67qbeqOlbfT4mYtt6s/oc3G5zORfN69ydV
+BFddb/mSuvMOYFOEH7ljrQqFQlIaqup54VlY3xgI3tQBjc4by0SkADOjeeLOO7i0Rq+uQZr8run
4x8OJEJ0MuK1kFY1PfrL3YoSGKva+IAwhjm+flwskEscf8hbeRoyTEFsbzTf1Se+7P1A/IMLMmsd
YtKLdrRlziEFrXSnlL9Gd0zNEVBucos3KtaRViHe4Lbtaq7wluLfkgEdR5yThOiYvdoGcrikm6C5
tZFRbtWMjbbdC7MC/0ugcZ2ieX48XZUfGi16Pj9WL/vETbmzMi1WDtRDeK1UNinRg5EosQuDHt/P
9gmwVd5ZdzpV6BpVT1rhg6QbmZIrLAyf0FIQMs4iW5+62sF0s1DtxB242J5HNeABd1urwiYh9Qbk
rEV+OOp7aYih/Zj3fGK2rExplf/JWAWGdjS9kMKRzGKlpX7eGlb9CemeRaaIZAez2vJK4ZRXi2tM
yr61fTuoconhalacq4pHR9wx54yDjt6gl2ZUUXwAu4zbn9VjTPjmvkaxLg4iHQ3NWUSTN4AZlIwk
5VvU9+Ym1GR6kFRyhEcTUvDs+X3PGYnuoL6wzRgJ9/8N1GoIav7srpkp2hMgJ5rqcg0MPB4evwFk
gFQLL5tMdIzvd7gOuRBSFP/EI3AcbecByy0ljdxFyHT7HMc0GlInHfWicshFtFja9zw3LoFTT1DY
VYo8rRsM7wvNHKDkq7kKa1ZVLCJMATMVyBldecldBXc86qgDmvmjwamILuVFKoUn71pxU02jFSu3
+p1NPQiNVE3mvoO259XB4gLIDK4nBuu9y//S0d8weRrVq7Ed6LcO3WT1Wya1Z6tam3+vmhdI9H5s
d8myuhHYFi9NMX1ZjM0/adOQELpu5Vc8LAgM3j7A8vyzLmmB46vFmSEqWA4KpJu2L8h6Ot72AwYc
kWIOrWLhc0kY6VOZnT0tcVQG/tQAiwzSzODV1VQ2kneMHv0DxGuofrHKRT5dsJItejdaL9jeJYab
6qpasG2JwcwOvq3WdbCezpUTuPZNFdL0bPdZjR344ZUzeEVM0wxXA4G+VbgX2hgb18+EChF12d4c
RZiN5mKCec8RLo6xj4S+p+Q8wADYbv3w0dwG/jeugaDZZhs1GJfpHQEXkAh2fZ4VR5H0IuoKFtdR
krkVC8+gt6Zxrx09n1nv9/2NcuAGvobQjC0djKqoFsqCs11ppDYn5l6p9oQ280HMeEv5egECL5P5
N9o8TKAKKOtpzgW7ffRq83RM9oq3YBhcsdRFubvzsDUd9yzGDHQkU085YrUsNoB1jSLK4PmSvMua
1BM8L8HOc0pOX54Ds+GB5qUUSpgQY1jEQJtukuw7oPfr4UdhwO35tvVIbDC4qHFT/Qu4+T7CGQ0p
5WEcRbWj4MypNoWObmsKsmtFnJpFKrBFZGZFVMdIJz+xZKFqy/q1jDnim5o5fKFvSNQVF2/G5hBL
iehQzfVPatHh2TK1KxEx8JIRxsoOKgM9pOHG3OGt30HdsOiXmXffY0GD+gMZaQWTbdzPv8WIfeWk
bJUFXyt/+25ke+CwaKlWFNZ6V8PSyj3HiVSOakn9OWg7zEnBn6jmnD/A+gtyXDORZAnifluQawM+
2eWyqQTrELeH7OtygZPNQdnYxzfpyEktrZgN7NEHz+/JL4oQu3OLSQHO3s7UkqRVgX8exlaFWUnW
rsodVNAd32J003YZolHDWlvrMcrsVFqwFIv/b77clqlIfHMNz1dFO5SFxo1dAACAv/mwWYG7M7qW
ROgo7wsPaT9GOtxSPYRcMLL1m+EalT4kvrnsjJ42a2el57f6IEsYS/bHajZ+asr4EBy/A7v38gx7
dPkfdYMK8qfkCt5umkIccylwpPs7p63bJjWT1tIm9RR8lnT/9gFict1c+Y8yUUhb8tDDBsCll/GX
qLQH25iexgWDwETyjvQkBSUEgu92uVNbuOvu3sQfLJ3W6F/w+rT8dH4D2EM0nffBC2YHje8mETXV
MzOtdNxh3WuAzraUE4z7c4pAMi89uwrtlkAimnFKAQJWhlUc36/1ItMACNor+nUWg9kMUnoLy1uc
KIynNCLLfHnu3UuQYRL0ljZutbAq2fXBMb+OGTHY1SqYc35VpXYSZWHYy404OHJih6Pgu5AFH4zZ
65id24e9DN1I17jYHxan3XQCENrLSzkjY1EIYAmDJ1KV2KMlBKu0PG63ItBdovwyD6FpLlYe9P7c
xFGO3HN6LpyTQa/EeGSDF2xxwZio6lvLqqNjAP63RWa58Kva/RJLqaLez4FqFdMKeO7pgaD/9KAE
gf5AEa7y1zd+sLt8rsXPJdlLfE1yIoq7RiYZ1V8WUhs9ZMzbP8PHO1HVVbpbu34wAcOnlnf+C5tr
fNfm9gV4bwGQ9dsQOi4HAxLV5zC009IEWQkeNX4jQwMZiOmRgfzrYmOhXteeF49JYa535hg1Ebvw
teRz7zfdA+gdTDyW/I56N3/jHZU8SsdMi9N/8DJwo6fZpkFiHH3YgBQDx4E5jt5cqOxc+Okqni+W
VQgnBwe2DQKrn3jD0kkz3i8Xp8nbyVC535lf9oPVB9Vs41A2FAu08JioPFp1MPK5vISjOjwK2O57
P0FGdDWdGAYSt1r4cD46oVGMYTTeppxDGifurSXHBnAMJPZSYNMK0i0g6LOB1i30CrriI84WScd2
v4mAGDFcOV1gFeAVZHspbs9Agm2+4d1RDbWUv1rQ11ORlO6gsDmo8gM+yn+1nXVjOTNFyeCFOdwB
AxxkX/7cvpelD6c5ueQAvaUTPsVdIuow9p4U6EO1zjPtS2FJoBMq5bS4uuspgnGSBQKfj9fbAtGv
w8qS20C0blshjxXME+hVDzX+6Fj52Ay5l50IZ5DwIKLv+ryyLfdRPtJwx/M3b3ANjC2VWXPcu723
n1IaNxyr1N1X0VPRVP6oXkZY+6X9bBOuDbVzhCVRDw/2cCkfdCN0CfO1dNEW0FwvSCR8vwT0xJY3
b2rUROgyFev/3aiPkwtcgSyhIBhW9D8Rf6GUZ6ZmGXIRJQ8Ea+IycgxKcJSJyHvpLfjrvAnTWt0/
0yS/jwZmOEagPJJztiW+ThzDZBUrxmTmcEF1yZj5M7XUWpHkG3/A8xnqQWBiCtlVDjtldG1J81qr
f5tUmwRyX8KXT6xn3tlfhsN/PqQUWuUiFIkIKPmkRxlRodf9rBYY+x9I57fohrvV6b6vvp9C+Ul9
hmEB3snhCJ3Wv8JPEQXae545FKVGfG+1GwVnUVuJjAOJHPcVPKrhUjnPNf/WsfXsDNszPkcOBEZx
Ae8+Bdb7VtWnBmZ+djSWdtOO9fU31vJzBtwRJb0rDCK0H8+4RPajAfsKy/6ZdUT9N+HYHzCBkHuy
KBuvw0/roCu5+Yh/yC/E9ZUxJ9gn5o3kkGBCO+VizE6kzbpSfpDFYo4/8sdt6g7waHlQvCApzUJV
kV0ml7H7AhqPqgXkFbgn0Fhjml8/JOP8R62x/ZkpnBEL3KGcU9zR53eGu93rERXq1kPBSmuAdO3/
gmENwT+1rdKICCQnLwjI4BcyaMaW6qy9yikaaULAEXNnPGLbfqvohcfDemSnCtIGXMzhPHEgmD5F
MR/hF5ScmK9LTgovIlVf9enBKEl64zByjgGbHFSlqDg7/xIco5Vnl8zwq8cfkLOkVXKNOFiD9KgE
8Uy6oqnFyk0PQoRTmJIyRfQ0wufTCv26+UCFMsRKlRNlXj68HM4hcrXpQRZh57KUWoiXrAVGtCP8
NJcUPw7r40JB1ba+u95ZeErir76Y9vpTIVtyVnwyNse2ZE2SZpzu/Hyj4fsth54a6RV4uHSdiIWg
MR6DJKnvFUVJiYliNPZwX2Q6Wh8kZGY0OEp2iNLWQ26T5Fu3bJ6lluUz9+x/oxylRgkKuB9j8yRh
VMjQd/vYrTHV1660hbZmZwUtHtmr0JICSJi6TNsXoy5spTwEFvU72BDX26QDWZ77c4rpH9eeZK73
QtLB3XaG6TvQwnthVZBWFT0hdQqYkiWWzdz+8uMTsePu9nFn/auIcy+WD8jHasCppydOrhUh7G45
XGxCJ5iKSJbeHEvvZ7m6IFjdP9X3XnxcVE/0ckdyavGlLYAl+VrgCLI/x/nFs/TgSEGQ4ged5oSY
3iZlzEXmVX2HR5q2jX0BeeaGlTk8oBAKsrgP+rgKwUEvS1zlDantUZvoOnQnQYcxBtVR2oJEGz8w
dgXA+Q4nXwz9zw0TWh6WUDtIFy+N2dRs+wMuRbrIvB/myMvV9+6mmeleA6D9SIGk8DKxSBMJADvq
K8jKiZ32vrmYE6x7gRzUdRJ3SsN1/2bQ8mQMXjQ/K8ruc3ZKNoCJB03oekUS2LGSHWF6AgEz19Yn
276z8u2fQFamr4kOyxotWUIFtEfgIgU6T5FT62njBy1F51ltCGzyVhmd82cctz/I9aYOjwnG9wko
/2IZRBlSWjUeda+5zuhk3323OrKxbwObsj6qzHcnQD194OlJpjcCU5JXA7G6HCF9560MPKmAVPol
qqR+iq3JjrtEcZ/ISrSGJGZeZK3nn4aRLdDr8IXpMqxMcsC+trGkjQnX3/1IXwS6NS3+lHuQa1d1
cU3HoDxRRlsFzhw2Dqmv94WCiPbWPfeYHRsuuk7zVRNWzpvgTBkDenJHzOowKdwBG6RuOwrCSDob
Ky4gWRAUSOFGX//ak50L8Pl774KuNA6O8kNijS98X/i+q7FTdL0YmclRdCQ6vPtHnAsMPns1RFLP
B7UK9pu3cFtxYIa40g9dmgykmm1TPj1ebPVJjJozAF8kObN9CiAspZSzEFp4RkVWAGwkU2eEA8jh
j+6Ptk9FogXiylEqHdeoIKhXrBU//eK5oA1hzYgVEoVcw87a4hNNFn71J3RHMXLv9hTLkkJQgRz4
SnP+SK96OIKImMwY6poTdlWF7PXzVUKXUGXW5ZtEJP459tXaTLRKnINHGYlhILJ5E3xSENYEGDEd
hFGeHXQw4kJV0hgjQHDqRS0FEGfl4DfBpmqISTiX+vdJ58oGbVL7A2WaP7mwmlNFWL2NlqVAt3PP
ukXFswwBFuQj4gfOoAjno4DfjofQjGbuZvqZSG9FrHoonqYWvhPWbXZ9aA+OlYUGHD5TIE+UM6g2
aB4DzcnidU8npcW9Ij99IYEwH6qUJWRDLJjTzfIb91Z6akIuToc/zVaNYImrLpCj2Dlnr0yQilj5
MVHNja6NbefzeXMSBBj6rthdKvbv9hk58ymEsu+H2HNATWX2XI4XOXmDlvFm7r+AIBJxaCBFyYcd
DSe0EkOlLxUWQtfclpUAnnmIaMbSe2hd+Kz+jKBFpnoAgXqw+IWXvurX2/wCPG+gI3futyl/kJiD
HEwTGGRmYde8rIqWo8wPjwYKJRNKJNxnU5b88Cib/E7YBg3B419NgJtIaXnxfEE88cW7c7FxVZhF
8dYgL68qcnioMUy7RSz/BsGs0stQbeopn9z/6dkhLRCiEz0sBNx6HMNZ9ZOJQvX5Kn2NLkrlGKkj
EM01CibPwiuKoaNwGs9FOh3axVD8zAqwh6E9l8ZlEv+jYE5xG4aCFb8y6rCja6b/uPqOv6giX6an
kFa1sdLwCBQAqUIdTPKpCegRapMi2b7t4ZOVHx2Ktq5JT4M11ew3tSxhPrYl6jP1bB5B5/FBW42o
xr0R04DtvE27uGwcDaRCKquTcLIEvIyLQnJnF5SucxqKzI3aCVlD5G/d/nuP06B32p7SseIAr8+t
cg+pcXkYiw0CA91ygM/kD5Q5uey1Q1DVHz0o3O/CoUN0kbg8jHB2BBI3Bo8WXzsLTVp6b/+FNV1C
t9tk+2hKokA3N4QWjRuRWkCRYAl8j582lJrgJB+zOvwBLIj2hZ4UAG5mjNzzWyvyVXsRGxcF2S/n
7+UTC9yTuvN9hmSCUaQT90c7ErNLR9JeeQ00fztSUTXLQqxopTJg5GZbax4HlS2RR93o5rIx1k/f
dWyByLrcgYHt06QQu3D7qhei8A73MwTSFiLqF7Rp9tFvE+Ly77XGD6RktHfE0eHjatYsAnB8BOHQ
MsVxhdJwD4IPym6QPWAfDYMFoqHu78Gv7QgNu3w3vZp9ymHBja7tl6z7nKY3PnrksRDDMoRj0Tg4
HSglRIVys6uwVtUpmNvNNyOCAV9uNimDPdDO3QulsQiWS6vHCZTQuKnsvjYKo2ONQVRmU1TNu1Rn
y8ub3eGhWssIYHDuesuZASHRVtzFm1kG6C4WsywdeLNzZexGTTdqd2hQ1yQPI4aGpUw1bTQE95aq
Xq7QyLEqL4PVYRYFL8vuDs4kE/qNav48zMBvfhdeEJBrxPAt7FO/fZv3JAhcLJNIwGbXWbyQo7hr
qha3VTffKCJBS/A42jyGNFx1OerHKJZEdioBKSEL7YDl3iSpYzvrNvfKu9WjEWB/MjE9MRBFFeBA
bIr0DEGVwyxe+Mej4x38MQTtnetTlb5oYISErh0emT3lhZwIhZuI40vMB+ogaVb9U1WcM0Av79IQ
3Qq80WEHVr5RinWoIfuQDA5L9e6uXsCRUKSUCZwCy09Cr9Tpr+sJnVnI0ME42QQEfCcF6+5dPxA3
iInirjYPUnQMgOzDzQqbzGJdDejVCz+a5dbWtDmPVVJNJSfM3S90SL3wnCKo4YYbqSoZJtph2TmF
R5Y1957RuGyx6n4+4rlZnFr+XKBJwx279i4ASKP6UX9yaQ0B61ckVYMkpirAZFAeLYRxvu54bxqj
pZgKB/uOd+wzcl244q55mLTlDRzhUvYsrOmidlIUBWMjI8dCppjic5PQgas9kyQMhIM11/KRz9eS
O9/OFW7Z9qpx0+Hgl6fWYaDCvhYkYEn5uSyOqeTZdvyGQHes3qA/hAWp3io8YddrEf29viDT+Bwm
yItTt3oVUDRQCXpW2nh10N5d0JNmRG2PhHX10k2kWRqIa3OlccJwQAYV2FLP+tyPLyGI+W5BnovJ
weYsuQ0fCeqWTAZs/1elaV9V2Wzjhmpkw49Gp6oUGJQ+jMEPJqAogeZEHhwqdMye7Wm+0Hx6xhmI
TIgIg/iKydq76kzmGtdavFXX1HSLA+6P2BBwcqOIPLYOMYdhI2/eS7d0XSl1TTYCND8cS+RuX/vr
aZEzZNXQQ6jH+tj/0IowaHhiFI8nlJ+v+9ypZ2jA9teiI//kWAfZAmEOlXiFzEL1jetakDht9GZz
9Y7gmCWpdeLmWD7sxvyPxxjRzEupV0VMKaN2UunmdlzhBAuSOYqmwOVJue9TYfYD7D++Y7vfBKAs
i1dstyayrPlJb0+QCWhxfv0kCe2lFlAa/FivEt2yVNs7A9z0QSJjYHmBIfPSpJaAI0K1l3Hb2Pd4
MA+1f1Z3MSZKX1cZrUekgfWusnh3N0a45nwjgNMvHJNq6ZHMrCVGHfix8hHMWdIvxLkojhkeOaSV
KNMLCoJhspo0aFZTCkwxjOIbsb3AOf2NHTA2gFEb7Xu/PPk5WdjMDv6r7Awyob3UNG0YBcQmXct8
0ckz5sGdOJxvEwCiTUOHOnIMtv62RZROwU8u+Wn64RbV4kV1QrKxEWKn4Gkct/hvP57t+oG6DJ86
Eqs2tZb0HgcL1V+kLFPhBC8zMXso3+IfS3CiEMskwpF15Pc+nFguYHHogeGCTYl3LkV+RwDmUrut
UKgn7JeUACw8/uJ1MQnFM2y2mMIFSh/jf0GEC3tx3asdzhbyGLdmrmGYIEHlvkrd2UwsNX6qvc6k
GLQSsphYEgfNy1UpVIyyBAFDTihOLzvJ+qondU9lT/gjdtSH/tq97f1AYG7kzqD6lH9ATP9l7441
aG9Kkhv7Puu998nVXR1nY6Y6QQPvkk8FFfWChYULbOdkFErk8a4jFgXcFemaYUZq3pNy70/WrPyZ
2ih1g0xo6Hxr3bWqHWxyz5ed3LCMgefAA+m//nhgAwkXEl8ObBaW7t907fdtKhDnzH8cLihXZ5KZ
jKMM1Tp4PQMG7ycE4aKi9cGMb291df66B7pdrUQ80ZFwSCr8s/ZuMaqZlStqmLkHWTryoC4A59QZ
ivHr6JmPMsMgUwVsXCh2IT2ezppgQDBe1t1Mw/yqQk3EFFHtOzwHAyHuRo9KxwhR8nTC2xu/MTAj
fvEX3h7BMmvqs0ipPcmOENFI8tW7g6TYBNzkXjhKgqN/Oy9thaqojXGmllzQMAm0lpYBk7cZwcfJ
mOx0C8Mt88YDypLZO82cnE5jvfzo20qLZpU900u2/RoromW0Jix4jaIAQ5BVDPwLMOpvyWFxggY7
fQWf8zIgsebsS1ARfcWQLwGmysPUlYo8w1FaEQHu49BFv9NNXqFe5C9WCNmb+NjBrfSLYyZMATuW
cyJ9ZWgoAMN/0X3hAfsjPEYwERrg7UPSZddpRIrpzaBCUV6VQClyD/St26egE23/OJzetv4QKZNY
v3nackzTuDvdjkdmEimNM6g9l9VfbISCWVxY/l2+WEwtzpcI2CFIjyszV0gkXe5ZfDV28AbTml8Z
ZeD9tC3FpAsPVZfLQIq8L4ZirgYpUaqapRrJF8GA0zH/zCbfD5Dl5Ec0aVoBgTBpyZ8QLarTpmEs
ZF5EYwxURc/1tlrEI29gPM+7FEAjaHkVnBA1oeRipB4CDLvH5D/vZVrS+jjp+ZxEmgJpbHxkmrJ8
ysmIjnjUs2rg9bO2i6738hadMZX24EvvfB/egeBQBfS9J4lp8qbld1e8PNoZRqy4zLtjKTbz1e9P
Z3jChkR+l+fx6HPvlAaniHnBsa9o8gLnPkqOWQP0g4tC8LfvyJTFA3y/28dTYccf+rQ6sGL/qIhm
bQzNquad2emO82krAohJWP0OjjgYF26dUJq3Hqbdit2yZGxT9xd8Oajzoil7/ZYVWs2XVpPWUuFc
8LeX4L9wiC+PibLH3ueayY1UFuREJ4mitC3g06xvES/FgWluJuDEHXMNVRS3L7PjXg3b+Gzn2CpF
fwSE8chhsZ8R8l+taEkjh9tbDk1mcGx0NjRfwGJerTJnu/ylGdMFwq9+ur+uzTb9xLwc174R88Io
rgjp9X+vmFCIp0W1qwZAvMDGsqTKSbT5ObTw2lAkiJ/2Lbi0ZbicuQ/DPjsCfPHXgQI+z6y3eptG
77BO5x+0KSVP3XqXVH7kHN4yAuT3PiJ2/b5/CTYqdkTlCRL1ItZDX6VGHqaPQfCZoxmGvsDnAMvB
BozjKF9VnebI31uIrvoz7lDN8U2lT+Js4PKSWHQQ5VcMIy3TbtX97SiclWCRYSVmKlO6UNzdAzS5
Vl+4BjwGYIDgL8Iauex6jvZTkDyDeoaCjZ4z61EJ1HBzAjxCF3R6py6AJX0JeBPUH4OjDR+IUGTv
M2bq5uB46jXL44EUPC5ZbOB0PVjK2w2mRsgEPIRicOuZmMVEUk1RIMuBertNOiJustHDH8fmZu1y
enPYaG1VXmfnT/KuM2ahk/cflb9+N1M8o8joAvrdAoFUQj3xB+LkreWwpEntr6Leu8HqQmmxQMUB
sqNZBcAZ+sG7/29Bmt9Tzf0MLJXaO4cWhFOXX6kX23aQbJjZlin1RjFw8pGYEVcCvicy2htK7Qu7
Rcz7lKjLFUoxknL0HHkfVclVZz0UrQMsiAMkYgu2EL7lOywvP3rfhUDWn/nYiz5IuK8MqpN0ujC/
ozA+afVfxu1pPzn7nUijqf/qFZiwQXOHum3XReOFK1pPgOwTxq5m0egMAs+fXq/lzkpOWdedqkW9
fWscREhwUoc8BV5if3bSX9xaZl47EJcvi3Jln7R4W6hgsTZagcgUA0yCuqTOEC0sCveZeS++mBda
MnfpIyz1+g0hGulSsw3cOeDqIAXjsOtV7MJbnqbcEIAdLc0ujJdrlcYbSmlPxrO3BRGXidHVC5eI
+XWa46sU7cG6Z+BZdh6sHUHSRoJCyXJDQ8v13+vjYXM3wOSGE/M/9ikWla9YoQ4gMaLsx7ApP+q9
4gxuvQxQJ0H9vmOjrJp+pVnOWHgrDSSGFXBxwDpdUXk4Qs/bvdcT6ljdoBXlLRzcqBZlW34ujCUX
LuSdPdzXP7KxgRK7Ea9t6xzW6zW1MAh+a4YtiQMltje2Fp/fouP6PxRVWs8B1mGePcOmjMxyO+r1
tqAEra/P8jkeRIuK+DqcLS89GlLDxCPBt6Pjut6BTKV5EVGSCo1SbljgsYgHvqsvf+5cDke5Tez7
5u5HCAFzR4oXgaW5/Q0gWEO51aLNoqEcbmkc2hvze6PycQYiP39FDbvprRz7sCLgdjpPpYWmTMap
sQT08i2BSZOerlTz8l8dGWJnlrNyqOeUEDWKG5WbQWZEoXhkIrv2ILL2wVhXK1CsDLOSyG5Nohg1
wOpq3uQj3Z7hNjfShcQEcYKW7MLr4/nxB2SOt8EH59SOWOm9Kzbbe/yFr/fu0gY8nyb2v11u4IMp
+2RS6OJimsrOyWgbRJQV3WGM/SCUIt99ENPd+V9dkvWdElfaQM2Sdbgdd9Jd6eM4mDC6glLxpTee
GTHGWquxq87PWi76eevAVXQFj+CQhRrxpl9/EOqKz/DBG8gEFb+WF0mTcp6J3A3/Luywv1ibZiBF
9Aw/fqjUWFNf6bAtlsotsV1CfSK+4T7A/hLvoltuUcZR8GKDgOzTzQeA1zJP84W+oCPvwCcGjZ/B
oAUb+3x5sUlNuZKQHlw/yy0lrKH39KBnCgLEuYSEOVPxvMRDJ5E3hWHo3pQInpPD0ceOLo6rYLBw
BGvQq8wcDzUXuHH+lPjPN4K+ahkwwRq/93BthyhQoN2cQa89rWwhDqQxd8aXkbzRtf1rn7FS9NT4
GZGBIfyvXYOfNd784nTSe1AkIQsWoO5cWGi3x9gVJvkjqRjaYCGxXgvLGVtQ7FmpwbGvJdCDi+dF
ow0C2dJZCY4oPTaUi/MygUMkO+0/VshBeHTnvAX8Wr2Ad3l3j2vYll3Nc3peT6jNftKSs30uqij+
WYvBYVBuzf/Y3J8njRN/6ZWNGAqEMf8Jnu1JDX/E8TZBuP58ZbzfSp509anxaOWEj5T3aMcjIo1D
FuaDP25pJk5EBiPR1gd0wAuW3tD9gq194ImD1Tw4nNFS+LUT00YKsu5bf1cJPya3PagshWhcKTfU
VA7rcg+Aaf1FHqvJd0QMVp/UpbzMDObqGHZI0FggyzpuKpLk0nxIRXEXV/V+QH+3AT92Q/0UHE2M
rGlO4R2iBmX6+X3NesDKJomUbVNRtg9LBRyoxm4a0IPcQefHMG0AApH+9KmepCB2dvtGjddoXFzr
znqjD7OZIpyKCnJGQJw0xnn6JZLzZGXFXaEWe9u7OLoxnpgsLoP0HPz9vwdjpn2np7aEJfBgDzjF
KQp5tL8Pp+RZ3SZTU+0n+DAsFxlh6fA9Mxnwv9zRcDEsc7bZ28TuVF4w8EyQpERFyc02Z9JEbY6g
Ft3nu0FbjbIBYYEY1QDjPpGycrEBoPjQQBg+u3wooQE55ihpyomTnO+NiZuvWQ36z5wF/a4hh/8W
HQ1x6ny+uYRmaOv0JXqyMhaZvM1CBm9Zetp9v72joJjnUkFBGYFjnk0f/btOUvL0hiqdrtxb81Ca
9fhFevjs1Ui+UnxON3Y6JacK0otSKxbSvMMWk6InCWz7GUR6ZDonUFDL589DizdnSvwlo3ufnm5x
lQIerZF2Z+aKxzma+PXy4WAxYMIwWz1YvNZSarBrwIg/ysYt5/MvdzpFZ/6TKfhHJ/s+zD05qplp
9ojjQqyIjeoD8ji6CS+ytAT6sBZJo+GrJnHGYxwkPp7ACan8+Uhc6KGKZn5hJ3G4oR/wTSpY+HTq
pmAIIZ6NURYU7feClxd9RGPYFRglweiR/umAkGGJD8jytPiaJEdPYkH+1wWRqyZOm80GT9TCaeiD
fMFkNh7QDewDdUfVUFiQ/7w04nlQ2w7M7g0VdhgCvpgFMxQ40nmjOPmNyD2gOmtUw9b3NW2JTm4k
FtIrYLxl6+kUdOU8UgC4wKyfJnpmM/ui3X0b2xden8DRN2AZhSqIHPO3Y5mcYo+xOi2bWNGuJoPj
rv7ZoFmvIqNsfFI0VyRHnuYzGowH9tUi9icEVu4WpNl2DSssXOJ7hQ2N4hvMIZ79nDxoOBx5rNFl
NY+53MgodUYWAJC6ZZ0IUmTcRdEol+2rypcGA6NSnFRbyBu9/B/TA8o2X59ibuarGLTOAdbV/W9t
EgDPLjPQ6mrjIcww+ysE1GAnC6T7kBaavCB3SKXpVOU5nRlr+3HW75pg5awDqFPzGPVGYuzrGzy9
7+izqREcg1fQAvQbibb2pXpM2DKZNmOSKc9gy7vRBx8iha7QDouUNncPR00p+Ce/yo4Cem+3WpgF
/U0lV4fEIxCEXklKAsBTeJ5d4JW6XGhqk6WgcahAGM6nhQ6i7d2YEWMw47UBCVTliZWNCGvq/mD5
p56Zpy10MlDEMs3V2QdBA5wc9eYtPCkXbup0RAQAGmxL+AGSDYAj+egzJ9cNjwzTjwccTnSt/OtL
tTxgVf1VSNFaYSeYEM6Ob9+YG1SMAEUoJkUxhM3JgmvWDUZe2ptwze1wLr73u+ulDN3VS6q+WHFI
fHOBDATqRCRvrA2o1mDVwX/RciQDHd6GhDjpIJ+Oi35eQ7IH+9Ki17322AlrdLFkgeKkQmFCkSVu
rWzxWVZGPfjcB++FhKfCQNMivcCSb6hGS8kZNFuzMKYQrnPxT2i1cuzjRnKTL325bDFIOaef7E27
JW0OjD+M+B3NyPv03SBuYiM+FWBUAHh8whERfW76nHm5GDX1DGgo2Pf01hS/VIpGx49T0X+Fp2Wf
zLXWHHqeg743ZN3693YUy57SzTSnP/E8H2gO3cGjl+z+u9Z6swEJjD9MOmBCg3/nmqX6neC3mk5M
l9Bi2LXdXHID6P0fayXLx6jf5eyosTkmuiMa3Tl19h+apiYRXL39jcMkLWKcgw8UmS6T5tkTPEjV
r1fJ7Ju0hCjS3Gsx+sVnMZAFmsXCfhmWUBRVHSRnWU537401RbtjpC4PVsbyjHXQjfpLM/ZYUlmm
0vX7zskkZzH3uN4xzeklSnsbxDBQefCLsQqLrfnx13/yHPuKWvI1Z5smMxPiagDo5MNXifuCKlKL
KDUAgbvdMzLv1es8Q5TxHtDjx3fmBbHP47aiTA1f7GD2HfXL8AVWJfLQ2F6/TBukn2RbuiPm7oP3
UjFzRjqsZ2Sdh/XHSV3f09kFcTlQ4NPrJgjk1k+MQck7tag00CyvxqwBh6cVsWBycRZKW8yGWjh2
UqYE5Rf/cxkTtbFQehs72dPBfMJGWSxf0CY+BE0glRbZhAFkZYLmlK70LWNMG2796q/u5gcHjcOL
YfwWOhqkgx1Fe/HOIvigX59QeyczDy0rGtEQmBp+mSj8MZMPxdQuBQHcqx/GSQfERIGWWncyVEOj
U0esby63aOw9jLbHWUoA5xy1zNcdQ9I/dHilX5A+9DYEgaKPJUnWOjew6Z5M8dCfC69bzWLsni79
7MblNd5ShsXbqf1NH51PC+BFKaRhlQ0edyVecxatCS21fXN2h/gBdb0UzoUQfF8dviNOrViFyUCA
VMlTo+W2JUlUrds+Ov3o8B+0nVDDfl2NSZuzWeGXhis00vmLbXk0wtvREUdXzB+iU5jGBy2tu+ZD
Cg+9HMx9CYA9hXy8VbE5QVjRtC8ARt1pQSUOoAlltABZmsSaunFIOFJuTlz491AOoQIWdSVPYG9W
MT2wQ6VB7g7fQEqZAnacmfVK9+xEG//7gJ1NrHt8M3XNBREqL17lA9YkEJsCuREoT4VnfB6xdzi+
W8Ku+ypRLFmgP7Ucjx/QzakzqTVnkh8BEszgqi5bmbvQtPPH7C1sdBy4f6UIbDAn//vS2Wj9F/O4
Li/GQSS+Al77cAWk75i8cuSF463eNGSr7VPw8yo4E9EYw9HL9QCLlymmC4xpMrnT9T3WmLBvgD4y
GkpdWN16Ig+2tad4zokRuEMCQvQPNISUB6dZEc4Wl5Wx6BwahJUdeKlHMPu7hD/Ay/JkVqNbXw4l
PisLfEtuHvlPGKsKZ/awkqrqGn1RWwTlEmI8u8WEDGlQsT3lTDhZXOJM3MFPomp8uv0GW1VjKodQ
VGBk0jlJL5BBlWTTFpoSPFSsQFeLfBecsOqKwCCqSw3w6u2xacogejlJVQ6xlw2VhONUMjvX/q89
dr/yJI5nt9aiEv97+Uq7BE5eA3Z2L3awW5DvzFUjj9aVfk4Rvlvy19kNMcNXDKQ96ouXXkTsL2B+
4qR/bfZrj2n7VlvQZhDgbSUMGCW6luZMYBFu5Ar3FCLkOLS5THOmfk3kvmsyF1oDgsrKFYdQvOgq
QLx3pbxeGm7USCkeFec0RodzFC/O761qK27dPOnL49BEUyNMXh/04/PmNAPccxTcfCvVETOJJTPP
BMwcHTVb6+pDnKtAVQJOa52yIWfOL9+6EfFAwPVNSwCQcyXOxZfJVFEIMrdTrHff2biKgbHj99D3
SNJkgbC3pmuR2YpZ+GatHl1L0TQy7DhE2urvrYZHlZKNLr+3aryWQKEb2wEZjRuttTY8y95b7xvo
+qsF3U9gIw/Wqof/rMzFt8CmTYgy2C4AWUlUsFxeipeKp+O2AiBBoI4J0bMuCXn/BIxMgjI1Mahu
fh+bKs6d21QuChdHBRvL1+t25RIwNisdSwA4iG9Yh/GeguqT0T6fY5qqyE0SsBOhkQmoCHQvzwrm
7JQIl9+f6PivMxbmgBfOrybvV2fb5JbM6ThemvoYJO8P/beJcSzmKtwBR2GTnC55H2Nx6s8+oks8
jzAPlKZ4chLgYTtfAhVw7ktkA59lzXJk+XN7LYuZ7jWQQ9hVqNCRt7C3clSZsq4LuS7cdDP8TRUb
FH8VbD7XB0Uen6AeFPRclSu4ScGrcpXVdHIbxUG38rTp14F4xvC9Ge4mhd6is4b23JPBQxo6RH27
zqGXNOwrSTGBifzP4muILo7Y5wjdejypb+916OW1SSbUygC0iY7PEwLciU4fVsk2vOfmFGsLoLGq
ExgYgMx06ToQilfuKc1XGUPdcuHEcQMqEvSKa0h1W8mYSqm13VXdW0kvcWkkg9jIk74GUccBG7hG
A8E3kzM4K5zplExuOBs8ZE0IK21LvJ/JMLrAiqEL6YESjyUIx04wxvFggOgUFtc2ACFVh19WgKoO
7HB1ze7H2wVzW22WV5U7twyyMJLf1VefLLQgM6NsJmrUFfq0NJdN512bonDxZB6lP2g6pVkRNa1k
9rFFWphooOshtnA8H+1w1nmOYWrcRT8cI5Vk3VqvG8YdQYGhq8vYo1BXl+F+bwVoaRavwugJml+n
FydZw7dOyiknAzc5FR3VbEEawvyYokU5AsXRQWYHA3/QR6c7hzmM5tu+c7FVgU3Ka9PM2EndXzwe
FDY8k0QAdTJc2sZb67+Df7F5aFLVW6octcO0u3hwZMbNRfB08eAZ/+wXSE219u8dGtHgAgR0mrZD
oDBjrWrm9vFdE+VYIIQzRszqzyWJVJ+9fY91RxvVi8qgcS501POMORi722Jn6QYRDqnbm9srwWQc
IWcqpgTsnxOTKvySqjysaHHLV3F+y1YFJCkLcCWynlWtI60eyUiKVsISulwRVtJvSSEzciEUlKS3
q7wlcLfnvHMkqtdWkGGrx1+WPzBObHpzRdQgVKcsT2irYrWBdx6YeszhsPQpUzLxEYA2w2+Dt7iy
bh6DHUpn40BMsx9xq23+kZjJsjG20FL9DQFApThVA51CZjOXuSzBfyc3g+FdNzKIKwAngT4FMGfn
0QqbN3pittbye6bXlZ4j7WsFAQnY7NmPTxcBhZV6Vz9d/2WM9pUMTYjuGnvr8LjMSGrlG712jtgP
RfbjFQpcwhdk4IMBTiNuqYQU/9qYeI1EVPm7Y59is64IiBId2LPiGF3998o79/D5zzfs6sDSGcPO
NhyeRmPYobaZXxURwNkXOop0NwkIY6/bObUnm5GqK5aL2s9WRKBYNyIpeGoG2hhR8wdUhtYiIoL/
jAfa+z5AD/ZR62efIhym/V/mAGVphxId1SbWotLcwU6gxb0QrNrkCST970O6nqcBSy6zi65nO8/Y
UVXtj+8450S1Mc0FZskhDNzBTV1sw0axmpHoz8kDCJJ/g3SUaVR7z2JersOcih6VbME+bN8Qle9A
YiZ6ovJnRdHztSVnL1E6Sju32CrzGNCdErA/EFgr14J1Cu28b3//WV2L/fpQI3EPoqzJPq9XKtRV
thQImiXRdqccvuCTM14pvOTHRDz+MF6z7QVEbJSjGu9vx2e70C9hqmKfXOmUazmcNT9o+rYhowG1
4QEYrnsUbWEffkoBZPuvDDrzQ3DsY3TsxhvDm8527NHIZkJjydqBygsRrgKPY/BlebrYnFMSv4Ix
6Bzr9N4fU7RH4BlZpJwru+qKbPz03Jthety8strN6PS50gVm3Rhu4qxouOBNqX8j3Z/54yJ36Eec
vJl3CnJ2EjdN0BaYyOItzZAUjCszz8T+zvvlq2ac0YK9cZxD3Vstv3JMEjAQtu6qCUKNNR84cnsq
318zb1QWfrxcf2LMHZj9nLOnwU/Segk2WfZgpfUmwastpzDiu4JnWlEKjpsiqAVXgo6VBK4/ftQg
oGTRh+dWAzmEFk7Gd83xmUW2qJ5Z8YdwRZo7qDt1QtC7loY/fO8bUH145G+g1sPDEuhD+8tYHQwn
9FIFDkufEDKlpctzzS1WceMy+QH4Gq77n5dTjbDbeunVMB/MaAkTvXr+A/DdKHt0VXugMi+NmBm6
Ls5vN13gQzaWiKu9SsA0ha65WxLTnvcE/FYsX5obJts5ZffSimk47f+E4IKussCkLJE4NV3aagtj
MQKTFKhd0GGKXi3wzNngFtJb6qsCnm54H6xhuxtTZvDR/m3M8bI34SlCFEJvv2uu3REaD0q2AoRA
j4OcoCz4ksHuUGA6L/Fl9mq/eaKGC6E1pfzMor2v/Cze3VuMUSpww7geYiTPq+VtO9GjcNBxZNEO
Jcu1WeGWrk4PWBJ43TcsVfKlHYZrA7svYiXnIxMtx3x17VzVba7RFK5YYdYCDzvhirnybvdN6EvE
96Zg6CXfGohPD0UY88fOZ9zYs75IeKqwlF2CAFTwW1wv5f/UmWo2i5lv0E00ivW7NBqYLMQotjBv
Ee5tbpT7daUzNEGtLpeuPDLmRQqlGZGuuSIBps9FCqrJm2pznhCXwgtHykUKGmmqk23Gh1qw3ZsX
QDxqBg6ZgwF+HfDhhSRO+9UPsY4+iLoC5g+GQGrO8wyRFQSuT9ffkJrb6gYy0m2IRdhpxjgGCToX
vhlffq4FYVfhv1Om/h3oX6gLy8I08sLqflx+khwUVlDS4U+N+9wzTpVTdmja3t1maRIbFGv95/BK
Fs1wdcx7OgJYiLL3tDDA6N7SGPieV1PPIj2uRtoU1aLa7T8oHu2D329mxMNaWooFuyBkEJ25lgpA
eUUDXn7wrMNt0IhFcnE4+luMSx9567IjSLKxvFAboS3PSCeYr4vmDb31/nDnoGECfojIw+8ivRKF
DiumyRs9mC1RiqWvbmdTk6wStRuXaDeimVA53QG6g6CZ3aMxyeGIKrf+mfSQV8NVMaelO7ICgPIu
6qnwTNFeWeIx87gc7+ZY5Bc8xGQHvhJJn2QptQVt+p5eD6TPfZdAq8o2J552U1mSiZ4ia+nOJGy5
QMjBJPbFJzk2Aage5IkKsWOUkLZEbnRsrERkEW5XJnvFfvHnyfMpXDnpzxnrXPan4o9ow/QSLSEN
8bceSHglSm+DGhdR5fNjz640ZkED1YWrtABzLD4YXjb9faRQaXV7VN1ogpOL9uKMXyV21oWl/JED
7kNetC1J8a3mmAMxLTRty+hbE2Xn07jEF/HkQgxdoSQVuF89ZTwqDeASF5IoqjrEeLgT7eiUO6j1
hbCVAxVNBbSp+aKPW9jxStWwug9/FSU5bIn4rXjROJriSwsqA/SSSWKbJGH2yFQ8/1mbHRjmrjHd
xADQOxPyQXzqM0jZI5uwPaSkmLixS6iIgzi6V/WNVYFiXQNviHNOvLfEF0e46O4U3mcju/EWyXMi
W3Uujv2s/Jjuc1nyAl9z48PhgH+LH33j0qA8eqSgj+JVagu7X1z8/rXSNAdKBL7PeZ7i7R0CDOpu
t7iOWnxluCggb7c3djI0Pj/NOfpK/beTro1gAn333PRJ+zoBP88KL1topY/cext5NUjpedCf9iTd
6BqZ3xdiXArF7f1MLAZbXWP8Lyy6hbIuyucHr/WRLGZKpuqdeUD+yBJJuLwdic8rD2yanNMSimHW
PLUk1ZzDw3Vyhck46tbZ/4MVBqidr5m0zmvxN/RoAp8kMzXu1sU9pTdXmEkzbwvrIWzf82uoI/kw
kO1wDNRrBfK0S2mHDfKvNrbJlUT2NUs41/e+a0a7gy1GQ8RCrC6Vrw9zXJTcg+8yg6Y8UPEIMZAY
bqV+oTJoaV4w7GqLVcPQrlyw0GM+l4BlJh26Pr5sHQPi4o7rXuL8yqzTAyIdEE1z2qiXdd3ZDUJm
RuETtwdKZ4UP3qcyP1KDx20ThEG70wGHra2RpA7K7TAkuZ/6xGQeYsF30hiWwsQQUd6JxzOe2xTV
tIJf/HzmJLORYugGJtWsZqh++CPvUwFjXs8RcAGCyLZdvdjIxHzUYP1uVq8dZyH/NiMl9/1Vpmbw
P0iX7sxIA6eczhOYMpdy/dfwQJ0sNYjXEERTTqqHgNeHbykZgxKpf6FDtinbZUk9IuX6XeAa8Lmp
UPNrYZ/XpAcWmKmETNyjc+ZmT2ttlUYPnu5n/PqRC6fq7y4kRq/dpcYPBeJdzSfsJ9Ct3cMe3sh1
1QZ4QClKo09V1JBqyiOYP5nGB86DdvsbLGxduPWkmNazpgikqlQDxCCm6MzosEv3Ety6O7ljwvZK
SFq6sVbyNXs5kIL5Y5UGQJwSpf5bLLH37O8GuLaZfc8Z96EA+IdIJWo69546+4Ymp+cmEFLJJuv8
hI482wnWZ2qPa5YVTyeLfZDVfac0hUruYBCj9hbIGdJ/nw9P9U/gZyAiFgfDqMZkw0P1KlkAzyuP
RLulFW8tehz3Ck/U7+0Y4kFODaUz/KxKJA6Zlh3JUnk0Lh27k+rFPwFy5V0IiCoLXKGsVb/D5Gs1
8jNd+stK2Nb+YMtSRGNYzlzRGIzF+8Ud1pf/WPmePZWi2iI+O34ybAhTGifUHRwAjg+kXgjf6K2H
i3mtejhYks3QcUwurerF45p7qiMgf+pHfW6f51+SXpd2q4wJ4AtxHxbdYKQ9ZuX6T9IAC/vGRcYe
/K9F7K262kv6MvUvbtgpquTh4cBK/yMovMvrU+up0WDgHkIDnu+htLoeT3PomsWSuXqrk23VB7SY
ZYb8fuiOVN055xVLICy5e+Hu5ZJHEI111gGgQz/e+zou3yNQJjxwa6Gyk1FKCSsxOigTJ1SNozRc
kFvLcPjAqACAb0Mx3vNr2geRYYjXlZAVGy0ISE2NTAo2BWUSkKHUY6T5ijHDHUXMsi8O2fC45Boj
QIsRtnXKxejZQfD83xzKf2B4Jt5beUGBRYU4sBrDNSDNoN5j9+4aaTybWeQymAAq7WHMWeurHL2X
hhPokdZdMucXJNEUgOO7sJfpGzJMrn544NxIEipED3q+ljBZIjLBXIXUZ0fddp1LUvVXLDzGuvxt
aQwEijuOlgB7Txs5rWZoGzIy4EPpYhY5IzleQoqEttjmn3kb/j55FziDCsydNsf0E5KAOrcqyONI
r4D41F46HftRTLk7+wEeSQomjQ6PDckB0q75c4qnHVv1qrVMASK9qJ43zB+huDkJCdFjpEY9AqXM
PN12aPkeDnFPf8d3WJN4TDnQzoDuGMASTNt/VkOhlgUswQ0hOK2UA5WDNuOCqF2juQRGCxVtArjM
RynUKXE0V2VCM7Rjg0FAVJv1M/hFKvxTpwmr6kjk6/dbwk1vwMkeJizdIoxrDcUJpu2CGkprM59B
LNxMooBiGhfoKomhwjwwATSLU9EB76bdGMr/HXFwohjhOIGMgQt/a7vWLb/SLuhLhEaiSi+sii4M
6Iemd/cEHtqxW8EOiBiTICTY70m9kXd9FAuMb6omHoY+i1NJea3lNGbmNH7JvMbwjq9TEkjjNWme
JMODn04AUBmw74iEumgfK/nqtb2v0ZP/5SPeuBRSJfp+FGuwgOh8D+kS33ViwpIjMGpxl90O3qOL
D82C+LOVbt5+LZf4auKwAwL/JbgsqWHrc01mWr9b4MNg4Sf8PiOeU09Wccuf/vLsyzoBQlx5DqY+
3IfzsV9ihMLOZ68SW3UjjUBtiY9zlFZfyejfPh5UCAY/OPVWvinHR8B8ZFNfMIEOfGcKgVcKLT4V
hDBwBmCW+xM3KNTJFEOcOh6/FyJBq9vMXVWurnc+ISZV+oGbQLkwsiGT/BQFcO24tuQEGqCmLre2
STFqlm3bTQIFvAQSRfUZBOwdPBpdMXNbW0Z6V59IJq0zj7tJvP6JfjvoeJOW3AdZBqHIDoYBGog/
L7rsEVB80w5C+nq0JolXpk9+dlyorWpN+CVoFXytWVmhTp1620XrzdR16R7hRJwNL7xH8H7hbgfC
EWmQHkJH7eEvuP+Z4hZPr7KjFODAB2DkT6HyxDw69yXvEAbdshsOGgNKjMuu82l6qESWzjJ0pE2g
PZ2uxgQ0n5eFHGBc0nXVOSo6A5JthT8qQ6nK4XCVmUpVJ6amseYv9h+U7MXY9ErvMmghEFcthJN1
fZcxZAp6cS6AnXIU+tq2cPTjabPsgUcYPixpjzN0gKr7UzA9b1h8R6qSHdtjLn2LPjFLb/m5S0je
ojihU8Ye6nT3VbDQ9PUAFKzyQ1628XI5U0bB1Oev1th0KXLbDt2JiLPLR0BPBIN7kFSPA3AOolB1
+RKOiFpUX+HLEEBbEuXT0o84LoDucpApXaxXp47IB6LFaOg+gJCBsWfRrcL+alYQFzcpgVbqdRVl
PEM7ZWHiksWlpJYcQmHYm7zJFCnvOlFEUC91jDMcFDiSU6MWcZj/SaAV6QSJZrDdr5FBOZfCkfNv
nxbY4nXZy+IBADdhbhAS5hGq8FM8FQI6FhjnB7tlPq2w5sUmDDDAvudyr6UzrT25Wi0KKL/DTy3U
IyNInXcqVBYhOo2DbJXGfeg7yPTK3801nOoeZq4V1at7X7sNqjTgzmfgrOuTu3gQQgnEryP6+v6C
NR3gEW88S+wCg8BIYGt9VOTZ80GD+HZ6Pqw5AJr56SiNe1KekDXgvUZOyv9PNRg13L+hZZLs6dq2
o5I3EW3GzFHHG5vOmUL3uWaO5NCiShNWNy+IQ8rXxKYHP8Kmiuv3Cxbrc4sYAPoRVKwXey8VpRc5
UNqJYKKfTS2lXgKEmQPEfacKHhKL7k4CRPpddQICGcLchow4Ni6s6mm8z/ouin1lDLF2MU/HHnrm
auiWtWxYoX3Ee1DuunobeLsTMQelbygyR4lEY0Moz0GYBTsgr7EdMrYuXWG22FcvnS2nY4kSZJaZ
eVYXtdMwDtb7iDGcBSg+xaQCe425Q31C4GvlYzk5IZqA/1x/mCTF0ofFMqbhp+Fd8Eep4/lqdp5x
B0MLbTbkvMcXZwtocpLAVFIlRahvTAnhW/j8sQQvtm7yD2gHgVUBsMB3q/irFwY7q2iJPC8GEOGo
zCP01XCnicGBbjlM8WM8F+j24IIZ0DiG+7NEd3xCzf7Jv5PbqkeELXPRy6ItbOohpMR4vWqAlTWl
7xaQ7RKWZKwc2VIWYVj0MN2jVZmgb2Ing7FMXF9U9AajDUzqKwn5hp4rDeJi7t4ERbnxoxEPG49E
zgmvBQY+2yymHO4mkv6WjYZ1N2cxER+CGFTdBQMkL5ZId9MpvV6Y6ZOOiGbPRAMwY8LsT3f9YpPw
z0WQj/HhjDoHOcz3TBdjGeXXW/uantJGXd54DEt9eHkEhsbYozWCrnILLHhgENVGF/Yrt3iGZ7U1
PBKfoOOSuVp/MCXfIviUDXSLrlSiu2gtiNrMq74qVFjXV3p3UCSUWXSxK6yjlp2MuL80PMhfi7Gn
RCODaSnTjS/Dp3irCANCP6exrWlHA+jB8R2j5x6Fkb4MQU2mhwqCLfRWYUrTUvjnIFO8nymG656I
XRsDsDg4t33ZJUczGUjarRDDjJPH3XoYJYud82+/RqkP2Z5nGDqfgNS/QKz6BGRs1YJYWzEKz5/o
l6T1uyPuLXcz4m6wO5Q9La7u9bWVeGUIRPQUZ4JGkvWwcUAdVjmQSyjGuO9piMyJ4x+02Tt2kJAM
7FD1mm6UlmB7TuzhkOACRa4kYX/sbwwIAzplpMWq/FIOZ3SLcPgSVOgBDJN06b8My1OpkJQPp1QF
xn1awCGNgG2RRK6ZLBJmPD58HJtIYZJfjKmhOdQv7CIcAebpITJd+82q/5rbiqHXfbRdatvlo5Zn
iIkRJp0ub0utRwU+2j4a+UpPlmTF9mCxXpKNFi4iGlhu47cQ8MJI9+Ozx+M3hxlYGqyb+nMs5JXg
DPfFHyXibSiqKqDYpwd3qURzNjv6Lr+Mc4t7tVtxAvYlxEkVUtJVtmisc8hpOsbTaxrkwhjUYO2N
t2sEM/x4y6SISIKLhKiAZKjwgmNaXtVJJgGOhldy8A3lf6DTgz1+WEWWo2DYx8ius7+oQ4abiBr9
39Phiqg36LLUqiNXgggiA65O/bg6DBtUvB6sYXAg1mPTyuiPUM8n6DTTvlkRfHWjXBU8olystf1P
ytj9obq3lI1bJSE5XjRe2ob3cX9ybbTMk7GgVuJWsaYesAjMfoGHZlK8DkCqrRFuDXs32ul/Axpw
mFdKOz9HIedI+mhUQzwqThPgaAqkQ9+S2gkHrjRVFVOIUN/9VLjK9LceOABF2byEID07oxUeCwHb
bOBcCzaYfs5HeSXATpxYChg/FAEAMrZCuEJl0Lw6CMIODeWZssCUeZYnaA7gNeK9xZlwmf6aN/Mc
YBBZkglEr5DKMbAb0pDbHNYQFCSqzqW7QOFXgIqJq/YfBmEfk/ZKn8DcBR+ts1Z580ZcnOLrNDxS
819115qFanf/VAa2f4NoNOVOkhpfbmef2z22dysGNT+vKup9g9eDh0XtP0fVn/hslva1P5/WPrBV
pnIMDtvYIRfgJn/39n+bbTyvT8t4VdoUFQwYk6GIziulBYQ45P0U0I+g6+QyrPyciicR9DZPkLFU
q2Qu0/RCaPrf/2aVYqRd45oowleGulbmVCv20lb1PQBRQ/25DWL0mGbJVtOMosAhtGPJOackoXA6
QGIIYLasySHi/caicKgg1eZLlX/2AddViozGSs3A8FuC67p6A7PtdO29wUzDHMHC9Ff+N4jXp+uM
ZutGYKw5dMtlSTnD/UTtJsD3JJqysqXoFHE+YQFrZyqnq39y8n8Vh+xnR+1Ri1rMWHbiSewErjZ8
lpwvxOZNafcqoxFyfBQVa/U0R/KR6ceCznlYmTZsmVKLI85RngAPaEW/gqCdwr6IR57qgAU8FcCt
GUlbOK/UGOfXI+el9HsAfqclvw8uQVDmk2QfcBsClypMaMdIw64Of2IcNfCmLWJRiTXx/SgkMkKk
pualj9Pl3RppBg+qkgxPWnfiDNWyGOcZ5N09kEsFuxnu7sMXqNDNeR+b/l/aM4Xo2JCcABSqObdE
DTOuwDeswQpPcx5ei1BNcTKhADdjr+4t+p4+vUQDMS/fp4pDIib3zP4Qq6MRSTju7uKP+P6AWYS0
GV074fhW32bJJwCbS6BzG6eZPq+xoZeq/W2cXJaOxLV2AgngxcwfNP/U7ShGN95eigCkCdUxnhrp
uAHG6Iu78mBKLKUgP4w5t1vQeZMoXgX9cxvF2rbyjaF84P2CR+wGZ0E1PMBwsaH6WPKPhURYUoIS
mJfq2apmYejK6DACVKQaYocWKXr83sELWTDc0KIxIQ5wXzXQ7j1eoZykxJVJ/podxNZXCdm6XOpx
wxbXezsqUtr6qE98gqaYhpQTG+Z7ufVtNVG9o+DY18qJGXqaPLWfNYE0v+VWSqnhMFFqxzWK5laZ
R0NpwSIffe2Ccz5MbVBhBB3lMtsd6GNaOFNeyTHSK583HoWVmEjG7aFDmQhc9uoU92j0jSF76BCz
Nxfn0z+T1coYpyC3ndh9Ens+bsfBfLd3tTf5vT5TSjdKcB8IK8Yhvnyx+/FeMtKEu7I3GuT2S7e8
d5o7jQH9G38Xzh01XuE4/X3vsMfj3iymkQAntg1GqINcEo/Y+6okP/DTTLE2KW0CM3O+MtfdMCPo
2RDqoeh0qdAFxyZY3J2dBDlTzsQYP3iE5kus+8GYN+OKIdebYCTCbY4GelyaRjIalAml/KkFkS/B
4IcdT6vHrkkyVQr7Mh7Splr2qHHHKIFLGIHa9ABETOjpdKyOaL3SQ5HQ23Z6pNScUM7vdcYDJ0CT
t3Hblc9gESZF0+2qxKHm/UGXeDP0JwimySb6PNE5qzUl4/mEJLTqb8jg73OW8YZPPqi+VA9TUVq4
0SWdq22FBnAt1TVmcu3ywkh1+4fJLKAvCxU8jZt4C2AGr6VpCB0FwyBObORIj/GPDC5KpMpLYxwL
L/sMHXQjvKkXgozQaDT7vi+wpsTZ2/Bj1pOl29MW1Jh2Bfi7Oyjm358AOHysM51WmJj4rwztirDu
SMCMV19w1qXs8Q9/3MkaiJDwmeipfy8mwqKarR3765NpP9Wj6JTdtu7o8+XFyQ0q+OeClt2KOMfv
qE8gY86pOtHqC232PbqJ4rASSx6W+cTRznsGXYfQXgtFHA2jfIq1b5Gy/0XiQPIiEIGaPE0NrZlG
gvHhUBLYz3QahptdPwcChf3fgf5KxUWceTj4m5/cLVgC03a0vJTxn6u1YeXhOewF9zK7V2j8gmGP
jJxkumGGQldMnuMTes+P0aagqgoYbKMJ6SJ5qPcUkRY9nI2VGD9eFnx7t3mWiLkIhNopSKHU4ZkH
EtMWq3TrxPZ6+klwP6YPWEseYP3+AeJPwi2S+JTX5/3XRN6fIa8ttzTMeN6p8fG3h7kNqki3mb9M
CVZCwRHHTMLcyF23mtqAm+MuhemJF23DEgX2EX+aGKBjK3elrf1PHuuk82rwaX7sy7t/y04Pn7nR
YPQ3/335TIixY3Es753VGqwvoInrG6aqWEpbr4ZWqVxz8k+WCejsdn7BrN3BqqOPOFO4vW+KZWpN
SZG+YvYjTmTpNqUiy2Z5HMUkOJkEEFFIQzCGNa+jBBSCQ5YlujDmeBNjrxHI/rE7yD6+SwdY2jHS
m5S+dbQR9UnPRrVcbEqhTTyR1PtSul7HV55j282JFjgSKfHw8jGRlJoOsKCB8ahmTXNJCAbps/Ds
Gq3N2jVHuTa7LOP+VpaJFRi3EmtyJQBvXKZkn2PCRU3rsio2BLvOQA/Ku/aHTb0WoDzMYpEssYcy
q6Qfdqmc1TB7ZTjGnTf2SbN90fFPNA2ZUodlHOcmJbMOW6CXLzrEOjiuYUfR+EkN1DaLW8qe1DXL
VA8RElyGr0fAki5nGjnQH56KPeJlm++ZDUqfLjU/8awqv2IXNJbp4+Of6n3UjLCblvDtzd5dnpaG
kMDNMLh0W4sJzYoQlwSmgjZoH3elX1NOr6EiKRdmcvIoqy23kP3AtBzJ4PYhg+FCRiaBF1iN9/e8
REYTlHu+936Zth7tMRakRfz97aUMtbNH9WR7/D94tpqKPzukuyNwbGWnqjLx4pb9jBJvBCSj3AyE
S1XPF7BOA1x4jNUi9Tqar/uF2can4HvX6JCjueI8mQ+5u8llel0W9WKLZX4YLh8FCp795blAsZf/
OJRTgbwnzkNv8nvuhDzLW2LrQSMlHkL+ZCl2I8RHDpT8wG8VrVJOl2YEdI66CMUcpqLd+JjSSzim
dtOODrcCwluUXru1id5l7PbVfSvKlw+P9blyExdU/U9+CLdg9PvmCxn9CbjeOujxD3+Yj9J7NRKs
tBlWKvPSzl8fBNsNRbqcPB+NHFbs2l2tD0KZzBU6t/as01B3ALE8vfdZfxQgJfnMQfZO4YQb1Mxd
qhfPh243It8bVwfnWQNouBOOHGFVHYctvLg/Q2yzU+0AGDKZql/z6pUjKHL/dV1DDERr1fhMkWDR
XjOncT7zbALcL1lBlRN2xhOFa4MFQa4Zu3jPiHo57WY3lFEf8eb7g6awy0NdvS5PQBoStjy16p3o
11eFeLarKWQedSmvBI7xB3//rc/48ZaimJwkOZJqcB8XaBPnopMa21g27nH2ZF9EKlV8vc+3rlw0
5k0/CQF3WPahT3eqIb/1wO/1ky7QNRYo96bbxDyM6dbxW68htL5v8utrhWvs5INwquzrzUo2DeiF
R59Pljil7LRvfewwQ9jVQuBzfwDiw3nZsOJ8UPyA4m8cKr01YJdLcQwMM9/Jt19Pq5BShO5KD89V
swX1HZvyuF9gNsJOq87sdJAjzZvrwI6kF6lzTD6TNgLmM+Tf6xHzLI0e/UaJgqGCj48GWtKHHuJ7
TaS+dmc9dNgUpkD/lYtmm/hSXdHdqLVJp2VmFZtuvoDfsMSGPr32QZRCqahV4Gm/R6GotH9BlDJd
VtBRoUbJapNhP7uWBx/XYuuOLl0ZR58XCS8/lk0b+wWrzWnJV191unrFZom5Fkc6FRfgK7YTCboD
+NB/ZBZSEON1rfwDgzgL/anNLgVPlibWe6aineaCymMvA0bucZqkS7sndT+RuZr5MeLbdL+3SYgP
ssqKBOX5JFKoH1VUNvTwskWZNLtvbLaKVLkzOD4nIcHUu2+FGYbvAdPWGPjT1551OnkR9otj+KTz
Dr9mrIE8DN60JRlKXEYLfogOkDB5QUZilUaHD6AdumwPv2AU9oYKrKWcvBUThjD/I6HqPbBQH/MO
4cVAJi4KGjtXmk+NBPHNNjQ9lhTDYVVju/tZJM9sthP12yio9PH5ypP/V1sNpJWtL2Q+jts1E/2Q
J5PZu2cfTOPApOFkjmkkvAsLyJ5BC3AGgeWfDO7rVyXxsVjqvfknD1XlYf/vV2HN/AP6HDDsEdUb
2BPxx9oN5lVlQGC6PByqjKn098cLdzqJdVJWOFdyiQcMImYlmisz9MxGWOIQfKFRw4Fexp7ZvApG
JiXhyzVrsbF0M7vmCz9PZT12gG74GuH2EXtGjVhxUuBuDllVC049ix4TI2tXIBp0Tw7xi5E6yxvx
TjP+SMr3+qmJaCsC44y5qSTai9gYOMaBSTtUu2kyvPdRq5cAW0layA5Dj5/2WhTkoLYI1km49EL0
q27qsXLzUPGsYLCU9WMoRbm7kJ/uEW2eBbWePg/YZUcURS55kGi1S4rT8uSFo8rmxy/Hx7Us/SCq
gCTjsnrLNNvY63M0gvVLGyshKZ2a3y0xFN6E3NxAw5Q0/8x9aLksFZGXEVBEokhnignBGKOlmt7e
8sSaMKiescuFwvhS+ZjlzKqQbixberxE+5FODu9Gn3SNQIcAT/0hTF4FzWJ1kFoGiEih5ICz2W93
indeih3yRZd6jwHUGjUywyx3y2zU5FBaGts6TLndvLamhRVzTqnEyX6G0gk1GMJ8//gMRFfNxVYY
wdg4vmNQ1SCeqa11Qgw3Iv3Zu2/JcNMIZESMKzQrwBAeT04WPuf0nCn1zhJLrnVSWUZAry4xWy1h
rPjtLnQVoVKHNNQnf+Sr78zIPYmE89S/ODxJc7+YECAGCtN23CUhfLhomCnHNM50k6UbEyXQxGtg
/PFy/xK45ArxlrDvI3qKb9abYDJlrQtjGvXAx4idfsgRXzHc4hDuhCNkmAtAM9KP/2oQgwWl48wf
GIVoFiiLGleqbmEF1XAupMQT0sYjecCM6o8Aqbx5AlEy9Fnw6kdBoonBRa47yOXQBs8MLCScp4b1
QTJMxBYxY+YIHpOMBwvPBsdYO+c9L1Hh7PbgfjO/py6LhzXCJqsd+f5+WqaLe2qxVd8C2zVeZdDc
7mW+0Wy/xab+bn/8Oq+wylB1zFY1J4J7BSADZgEg0TYVYWMPBorOVeW2RFrWQzhCSGRkRRjX3CJ6
XVyYiosn7jBKzUbnC2PpoTQTmo6Zt/v4eehILm8t99ARzd3o+jj7F7zCqytunSmi08YEAi8KESh+
Rb9C9w9b/3Nj9V5OlxBYlmGlLj8aydXTp+Wcu8+dNT0bDr2+E9NMlJlTASxupA5fFK6MGrhrFjPP
6nrpkAHWo0YOKY29tk0+tkGjCJmZJUBPuAqu5gnLDuNXcQUfAs1kD7EURQopQI0Z+cGQHDm0FcU6
55gkMl+/mgG4Zq07CY2ktWBPytKyqVQfFnU33aJHkCX1WtvVM0acidVveYpGIgaL3IoCxGtV3Rk/
MT9p90wfFEh1k90lCqUiW5SQFEqiYFl5wXD3Wj9sO9c+CASUIOGEc7nPx4YbkKXWeKd3PJYWaodG
T3ag+KM7VEa+lW/4L2xdxVml0KLXQo4JCUxtbIdVWZeSMRsxUd741maeE0URYs7Y1BiuGGAxCkWz
K56ppxSV2DOlzCZhadeba5iRH2R+kumLD4irXc1lXBandeUqyySm0p04Sqk4lgISHB9IltICFFP3
YDLKmQ7/2AIl9lEGf+D5eoQlpbZvQ18giz47LMYsxOY1zY2UD0pW1qsnF+FFQ8PoHI6ZGZ2m6nuw
+gRDsU/VEuhLbwPEtvS7n5PdRsgsatl/AMYY2HCHgMmns6zpM4cL8wKck9DVfPnKjH1J73Fa92xK
5i7sILWcUK/M+Nw/GXQDxZCohIis73B9YbdiwLZGrScmLsuxJz9518rM7uOiF0+fSgGn5h6/9nY2
8ui7bjJ4ui+y67awo+NWwumpR93B/zWmMlC2VY3gBNlRSiV2gWREDbhA23/Fj/GxfA6J9zw/lnq6
l4vMmtMAVmjgaSI2HSiiqNNjP0dmzGBGvY2+AKg5AcxO5lZ9WpUjfyoHm8JQaQf2lWO4tRJFxIlP
3h7DnOC7EWqh0kTW12PA16cPPcOOwBbd1cM04OuQ0x9WfXrrsLpkirwb83H1ebW3vbcFwMaxPmgh
R00/N9SBVptwR0NuTTY4WxeiLpeM621/G5pT9ZoigVmxhnJ1AIxSyz4u0Z+crec5Ktw+7y37aotA
RWndpqXKEPHm3rKwTPVJuqzj9gEBiwmZmCFjd7DriZbqhjXyzvpnvvVkSWKJYKJLSLjnMKjFiJ4+
HbztNhNvrsB/yslncC2Hslx4ABs1e4ArwbzfRDadKGLmAN7gCFyIwO6axQjnon9R7UCmOdeZlbKY
FFjA/R9PCw9jxDBqbnz6JHqVXNx0K4ueTivgzv/vlaazIcUIDohNM4fv3Rzx2UkPgeFizqMyIVGp
zj5x9bPQX3GPujPdyUNIJH4y5GqiFrcQhlW9GSc5OU3w4FL2MSKv1fcM0dxSxusnijU5GwCaCLPo
00CVzNwgr1yjRheHYfcc/YlU+HaZiZztxQUbyfkMhhr+Na2R83YS/XnzguePvMnqWiyrUT4ULuSX
VRPWrcUw+Wk1QPVsCQyEslYKmDqbeSpzCGQ60PRMhlGAH4R1fxiVS5xUUgmxpIvxOWhfOHPOQLNm
p5aGr9VE38QJYs4BrkM53ivd04GpVNu5r1yHCMoVCymmWpV3qCKuMEqYwmdtGQov0HS7PpuaStfz
UwaTCdOyx88xiiC2eXuvf54+vOyjF6F/EmXYbcFwHXDTyEPd/IqpW5acLHG0zDSdS1Q9KYOp8ipk
jXwoZos/bkPaTbmJE5Fzq7fbFtV9aXDDdmBfHS4qumAWLtFSN/XtNRNrt58YMN8T0uIgssAoeMXb
W1zBfZsmIfcCM4MhCfUT7Qo94xHUotgmFk2/8wb/dT8evMCQUDNt3fkfH1y5DWjhpDLNt70BrdFY
c9AEmKSyoiTMZJdmnuJDLtoavJ/BBXZL0IffV42OpyG3AyTHJkD91nG4d9d0xqoaLGuXZr0jcoUA
tUe+3SdGYQFPwJVak99/CLI/bWHxqfdhpnAliecTFGn6cvhqKgvtYhAszql93JJ19ubH6bUjVu3j
CsKGfPksrh28PhwDP5Wq708CnC4ukEARpf+bj5D0Vk3jKC+TL1OGYysCS4vqLytcFem28TID6uSH
wAkCnSPqsd7IIKSxZnUH154SKrs9X8WE6vPDQoS8C0yNSeKsCiyVrg1tRCtIjGAUTgqyvHFVREjt
a3wATRyy8efr+R6NaUdf2iAdflos4UAb7Sav4K55ti4ats2/h9veO8bn2IC0VAEozhbwvAyVSFox
MTchdaghenbEToySZIVx89G9ZjMHOMeN1+44dGxN/trkz6zE5lVBuncGrOjGavGQbXck/KXDxqjE
l6KnZ3PxGLSp8W5y2N0v71QKMZTit1Trgpyh/2cYE4VJeaa/zSR9W0smMrm5bA+IhdIcQs2zKZPJ
7uOwcLmCp8LfEchjgpYP+S4dFHQZkK0/8we4PiDuQhiWBHsQqP8i9ensrFGoeoNKqYk17EbQo1rH
8bXJDxf0hqeYklt0acUaJ5tzWQ3Kr7EtHzi101ErZstbzXkG8R2KmuJi+2WIhDyK/+IviL8nM7Ib
3TEGBFLfNE97SrC/YqkNHPiRCHEM1QiRIgmk8QuHYjJnrasxLloVlxVt0ag+acEQ7OMRSRv9fX6B
Mk4A5h/Cf5rWSqKc4J1pPd7XvrMjo73n7tIKikWbkFbw6Uc/M08ZKvB60XlLC2Mexmf8fpzd/SCe
WgL4XvlALPouE9dhtFocMpMs3Fhn2PPB/A1tUIgmKZY8OkhecGj/ShoBSnP69gTXI/1V+UIJEUqz
H2KSRBzmywnlCj3fA7FqWjQN60WA0iO4UIrIC1FcfVCMSP/z9+U2zhUB1LnDWaB1M2KXTaqeE/RT
0cBaMQFwDXtuLmM6DMbDw3UxwWFMtg4gNaD9BCZUMlo/d0rldvYZwp7cIbiROHCs9oFolkFe7j5x
ZTkxqPdFROqFfzcjX/gd6JxrqzRsHgrHlzPMUtq5j359cBz1sO+Z/k7Cbc6Rf7tlmXlRkvYHpCBD
g1rp8LanAjZhdsUbeXKljklK/BSMda31Je7EZMzxj4+bqrpxHM+tWvRU481BQ1hsXdUBt4LNEB1Q
1+Ml442CWrLuLA9/bQ2JGD7nvIRDeiKmOr9Wmu8Cy94q8akuRDXTnPhK454MhPxsIhUOrMf/fLsc
0aMK4BfsWquuSfU/No3tD689VTXAygcFpFLM20npVe0qCtxcG/SKIwzmPVTi2vUYeYSAYnyghffk
5OKNSc2MWUrlwxbP8PCtM6WsuiOMs1KZ4SOfvh3DmwLmw3hP5bLfzvnop+mU6+FfFeWZxiYmE4xg
jcWUPd95Tk2uZy0sjUQfITo4dpzMiGE/PJlIr//38lTKsxXfR/pMxUlVoJVGEaNHBaW+u6lB3+0N
nlTPMUWueOrerQLQvm4XUdXEAQVTKSKXfgXDcvjIPREHvkGUYHvPhLYtmoQWGu5nBW/16rRANycQ
r2NqSyp+OzXpMFhS806CW17YoFAYXG8fF1MPwg7mYATRmEDuR3Uu6zdMKKWSOw/aPqFJ2JqB365b
vp1se33Lqy7bBmepKE90lV37l8KeaPB0j1DGtIMgaoN39yCTZyqxq747IT1Dfe3LiY7wufmGgiNx
Bc5PthmJGjGx1OQpEaIVAkwNySXjXnSD/YRKPCv2db2KICiXABJf3jiGarFOGZZEN9axwgqtrtVS
kVtrvLxlPH2T3nEv4zp5os07MqMCdLbvoC0YjCVvHuh13qe/RMw+A85RxFw26nroV/hddY9hmmP1
yHtizuyB4rmJCSW+O27X0JqCozvQQxHILYh/S9asU2q3sXcz8L9S9nO7g3TSNyRp3XBT0+FeWrFu
leIqdMymffvPNEYXodpOaORnSNLAji5QOoYnGpisoJNiuaxzsbeE4cYxzKkD3Vf8fOw9mTm4FtmK
oqSiaVF/edISKAgKKjvub+rL/fXtUaMvrfp4cVN/7MkEoCGJ5TsifEI7yp+SY5kaD+VS1Mha2U1b
qn+EeGSbAsaFf3LO1TVj0huFoVipFsK6yyJJ7+eSxCtw9VzmK1Z0YFWPT0h9zEUWDlu4thYGt76A
ScBtxH7Bzhle8f+A0I8dKiXs7K1rpsH8YZIu9iggULWbLELl3i9bSSrUviSTLjbCfZ35TfUM+uk2
zz/mUN3MMvX2dkCZO5jMcPlti+Z8z24AFDWfGFAE+d/3bVmqCqFjTYA0XsY2asZP5AgVM99uIckP
GUTP8pZ9Qc54GUaApJqMttJ+UXP6vlk9zbieKW0aCAZEI/OLZkx02UCD0LfBnGwgdkSMDRNgx1wt
wwXYRSYjjWIUerC4/10grQmWAbiTCobauaE7zGVjJKc9pZ9V3eRwWntoFcbrZBuyZWnofnli264R
ISkMhoy/5c8zSbvSZ37BMBN51/cbHHnDIcdBa7I1O2nxch5WC08xsnYMGqybBgmVmxDxfT3xuQKG
d+MBtI/Hp80MzaVb6cWzdAoz0fJy+eckg4282vLuxKAA8U/4jTzHzuIVYmJMjS/poekLsAVtBbZk
PLBt6GVNjUmiTfoAj4dvP7b+uikKB76kcEKaUrTzrynvWQmtW3dzuX2+JbPL0Of70BFk6FgUyWqJ
8vyMsL5IOKScEd59GmU1hLUjeOPLVP6BuLhkkkcQmjbz/o/v8Gdzna27EaA8oKbMQ78Szo1sczdD
rxgCO/WrQ9MaWTtcxuK9CPCktFBs2vDe/dGP/lCLQEAQEXCYE0EAIfTQtoXIWWEzlSJdeoHTBcWW
2msNvNjMEKSm6qSAlgIlUcDCPEu2p7ZRxEfd7xTccBNtDBfpeSxJMX/TFJQGdJr5jvA6ip5YLXGo
Uep7CKJHTgdsQUt1yDIWCYm1Iqlfd2P471uRcRQCMvXa9JB3qEZVY6OwTPK0G4B5WSTo3MgR7ky2
Q5tMQB2uIELbosJyKlmti2KMWFPYxBzvqxfzFZ1GSOp1vtfPsL37u0Jp2kZgaUUc7qYmUUIjG7jG
WhVzsxk7msVesKcbEBNoHJt3OYAzFToUyliazU1EzyLSuXBR7W9Bcrnjmsn3pPYPInVU+sgNYhPb
gZbqFqSl0WQZN56ceJYygjJcE0vd7YtD51XBtgl9y0UhZX1savwT70SnlAMjj4JBDYQXmeXyoR0I
ObVuQR39U2uyLfPTKMRTaaUfXxiVuPv7eder4XOMdRN3p+gAH0H6CVgknm3KeAkq1HxSDjVfwdCU
TvkM53wMzkUw8lKqmbNexqlLX4h7BuRni6sddG2f67AiAW6mm+m4q6RGCA0gQUjj9b9YYTFiUzr4
q130/NOURETTDlNubeR7xIgbSGJ7SEAoJRxQDJXZUnekFqziURNaZuKAKFDzsfn5PgOZ/9Wa5yBi
XAL/wkT8j+7H/Dn5Rc3KmXIMoyzUCS560J+ipLIwyaam8oHqZwIAHA6mD/h3pK4gBO3NFl39vwyS
BtBk/V8b3ehgflrAEZUUsHp9wDLtZ6wYQkaZriL89ZU1XNUtuH1+Msxb5fX2+66LO9+qH0532VUC
xfD7TT5F21ZdQkmhv7sfnVLU4FYp8u2Q0z/p4akGmCVfbgds6xExhwcwFQsPWsaygxPNEqgoKq42
0mxaw7uhziFa6CmrNdlHgcC5GDPkojU5jFMqZdEICpefNTAR+zI1s1rS25k70X9x/E44LMR74eI1
pcUXtbNzsvS5UvhNIIytEJ5Joy2P8QcOeTGsOy4pRVTtV4j4nR3TJWg/1MvP9gP1ttEypUfJy36M
jfOQ7Oc6E93OM4jnDus0wq0umLBzZe/2CKfXxthzcY97IQ8ya2tEqnyOoHIQct1kKfKdmrIPr7kK
w27HFDPmORf4WPbuJvJgiaoUxhWDCakUq7BE4werDYhB5yWlylfwl+VU0mt/37ehsLqNqSCJXOPj
PHkThkIGP3xLrk0uN/srpEZMRjZGPDZIUepTlKWp2LrRCJM3JzqNGE3dZi10tYMuYzuYBaM7LEgt
NR9hzE+lbDq7Ho+sBPRQ0Hc+9LBQLMyh2DT0NZVkUeK7035Kbe2K55GjkwC6RlcvXLLig4zDt2ma
mjrZyesznGDKayqvcDBkfL6RmJysQU+ErARbbq3wdccr8weFtiQEyynqqgUqRS4yS82iTPnSoldv
1bQW78gr/nPGYwga9xPj+NQ4YCZd+sWMTgaCsqE7DmkY4DC4bfeH8TsEFjDgF9hPSTt5QCBY4XZx
G7CbhDV7/Fx6FiTtGgZ1jLiI1fd5oFscj3UsTyAMr+MWRwShsYQ8tqEcaY35MgbDwlLyp4n5468c
AN3XFCax+zERj184ojueV2iAjmUEIWhVi7zGTVsDS1yBud7YFXWQQCcHLMf1KS9Do6QnYbqwQTSY
8qx+YzcPOJaZkr8oq5aekbu9EfraUeRCnCsFfzcVj7JOOU6pD0pp/nF22R5D3q/5H7z7RVjGKRsa
7RZZVsV8cE6IOi3HQgBDoi0A3CCEspD9l0vt2DACJf//YSdhEe17WPxmg1JqRVpac7Z+p2R1mvAn
rPYV9sxSEZcs7/vdB7W4yL2rOLWhc6c8O260Xkl4Zo190lIydVCoutHeS0eGuZbUDsMPF1kn5Y9Y
vL/d+GnMdfRD/d8ndOGIefIAi6Atqhc9EPLBuu87b2kahRDSFwPE7NystdNcsLMu/QtcG2SVZDFG
QMCrww0smM0a5pJg8xi3i/i/wU5PqUp0eWjjz+ORjkhnqJR5grbzWXMumX2EcVRPDLd9PRlUTNE7
OspnAwcoE9oDD3EotKiEt9cXaKdUEan3k6HHjaXu76VNpKQTeDoX294Xhb74IBDDPUntJ9d73zad
zFF8zXwfjfV9/Jr+CxfVKsFc4Xvk3Ts/jZDNsFJcLh0XnES1B2Fijv4aPJFhI71c7arMEhZG/cDv
Sue0LGLvP4NA1dD8vtPowkOefwOujAYwRYBb0/a6lJ6rQaXSzMOldsodbPnAa84KQb8CTwX8bBxX
b2GxWCPJkzzotNsnc6IsUoHvxQUFQIhEdJihPHA7T+ZRpIsAYrX3NtJMT9+EUL2vM990S0sY4y1v
AZ+g76tZro91VnqlgLuzaJy8EMyYlxyCrrWh7iR7ZPPueCqjHwchCehOcijQUPfKpfoBJyAG6Nt6
i7l+fI+yrjWzRluLnEMDI46FUQ95njZEzrAoGvgNv2c4fC29bGRoRTMQs9MBTA+TwlTyYMdePcg3
4mVExdezkeVFLrefLbxF7jV0QllnrMjGPRRwLrojLcoZqRlTYhEppjgohdFQ57NFI+LeS8o/GrXp
oNonEQYPxUGde1HsNK5qV2Bb4dwDsGX55BMe9yNfteRNMm1CkikuskCjEYbGkYrdKpTjGhH7kDcF
c9pFhm1gQix4pQkP6PWTwIlhAByDRfjOBvaTPk4th963/HRLCYqKSdG1shh51ic6gSve7OE18XNY
QB1eMQTQgfjlvf2IOZyceM2xa+euXStb48mfxtAmXk64YLpJiwf2ubElAJv/JrkE7UOoroiVxs0u
bDpdg1FaVDclej38IiLrvH+09pGTVqtZ1qiQsl9EJtyyr14u04CtDbaKxJ5oMgWRrMNm8H5AIrL9
j0fWOtUZ/RJGgGHMBhzcDqe4N3L7Kjq3glvkKARKE1TQ1GY7Ue9bIayx0Uzr3Jn1xewaWArR5mSk
RKEsER4nbhui4CEaMtxQOFt1axFf4XBvMSZHSJ8fq5pCKTI0W1MYUIdje6GMisYlC1kzHx6UdLhB
LzJta5MiiCmSAgHHW0SDjHa4iIGcFAYbS+A4usFpF7orc/UiIO11x6b03PBq46DFACp5lDs4Oc/e
Uq8h28eKQRB560taHMYxu7lMi2xmw4+HRNtGHovofepj+JOgsarcndFfAnUoMvmp7R0HrgjdbZAe
Hc9ue3D5hcyeIoYiuE6MhS+a9/sgrHr+IjjtsyxwUxA0Ws4OEOxky4gCKUTNxKnID1naqL7mJtbn
SQ8VdKkDs7ypJUzsWi9LonetoYNFxTyXsX5YlzJxdnxaa2vMbYTQkAxrEVqvyRgsd5bdMjRybQak
fcxsIn1lYg+HTm9839s3RsRjqCUl8Xpojlhe/Xv3hG33Y8mRVk4ZHGrkedBtuDJhDpRPAqK2Uupe
FklfNQfObADoCNOtXwB1ohIhFrKPKOTrMKTjZoIlGuqeWPIjpjG9gevAnCBV9yUQA/Etl67me8qB
OGWeQoE154KMxEQIJLKol79grw3BT7QhTPVXYEn0SqAEs8QqKuYveVCh99ep+VRZpLBFREonsAur
qIrzJ8+f4JD+2x4vv/rpZwyZLVciPAt3Qr3F5vDG8RbTlTXI6MkJ57sVFzcF4uFBiwdS/eZN/pxc
WUBCsKHJcL+ps5bLuy9Ffu58jd/WF5T8KZMnesWTvtdm6HK6ePZXhfhuGLOxSJujjY8H95s4zfAm
tJPpvmco66HVaEHLqwV1yNgZT/ZWJCYoUWJYOahlcDeMnwtDKXWnBIomJ/l4BsgmtsCujhY9J2Sj
VYpO5y7yQqyo0Eht1p573riXKptKeAF1XgSgerUVvbgVRkdlLs3SY6/UhliiM/gjgumeLRFz+xmr
YkTv9HzxLiwMqG6YzHQo+/4sWRWmnRA74VNQQDiANZfC5NL8UWUkBsc5PuU1pAm7SYlK7ggD1DFT
dpU6DRs9WtKQHCvNeoUUDu5AT+tI0gq+cRDK8IOAagMx2In4OT7ws8mLonQmaa07D6PwHPIFXO5J
n5Gt8jJQd5h2U23ulxOWbSansaC02efWMbrDaZRplAijvcNReaxeUudKjILx5Go5INUGhKM3HeT/
/nUNWY7mgbfyuAKgi7stNN174V4KELvRpf1+mCwppboittjYaUW7Ywv++6S9vo4GHh05hbu890OI
oemrIDsiYAOK49JfF0RgdnhtYBpywiNWB03nmtvwJjJphY9x84MFTa+4BFYJ5y+fvxmAHw2ANC23
95SMQ01Ciqf/y9FUd3sw9uQEBPiV3xbNGeAcVnjHKmAQrLroHzH447h0HeWYw+wqJLrt5BNln63R
qywdQ78Dx5s1jiWcevHqgOn02kfCHO3QJMNOuGOzy1LPWisX5sOifk6Ulx/e0APNpMPDecFeO1iy
mxrSAB3txX863Ea81e9oWu8dNzRrZUYYCCgwweEFazOW34C0R5QTZbM0j+bdOFz1K82cF8N9J/w/
/MClKPHvFwfw8DgyxajNZziDARghNt6SCgbsgOJN8Uj9PGL5mi75IKoNVB02kTbyHRPh7yVLi55q
T7PjQo8v+h0fUkFg4Bbc2L7fM9RIU1WKiPBk4dFmQuJ8dsuHedhoqBuSE1QFhZU+R1HB+qwTsC1M
LLtwRoNUAm39oFkdwvhqKomOK6MTSCfzR3KL/3FPZWZRZKXKEYJO18puE9DLpauA21RPHVzsDt7z
p3MB6JcTVWQk8vHrYu6aoFmuHc5Wksr5M1mYvIXwXvhWafsyzni68sxKXbgn6mhdH1wSXHgHJZ7/
nKEwInauChqJEvKD3dNFCxHuCeWTOGIDD5mhu7RtH1XW2NrAJXJjAzTqXs13BeAGT/iRrRuyKulT
rxvNjioaxvRaaI6k/sGF1WQHqEmDPUvsRo7xrnp48zTeo+0tuEtY20Bd/e4xR7koXiVM+sn6pL9E
rugGL3fCuOZ0aVackPdzOnO6T/rltttt+Q2eCV+3AmT7CFDCDwkSM343G9MD/g0lcAiGEZwBUES9
KTMSaFuV5d68hEU1mE1g2E+Vy8S8VKeOeQ67LkfDkpfOGdQkmexrSmC0KaP5g32RZvFeZ47BcljJ
JBHF/eS0tzPu/0ywOy6vUnA+7gC8vuFHpT9zaQlkp5Dn5i4nPlCOvDikNw6cvJgS6Ofq9QvLz/gN
Z2wxcpzj3UjuppM5sDmna7uiwHFOLLF/fTQIZNUGPzJPhEd97o9fxgtLpAOMmhHnTfL30NszFLie
8f7QUwzGTustoKpn28p+AHssPwoXY37uH/irLKz0eatQMNxxLL+pRAPj2QkHEA6HA76NqiwmI4ZK
2QnauJtgjD089cNelKOscMuoaPS/syuuSGhCr89euTq67MwtwTTu/jBucS5kyl5P1f2hBprvFBr1
O704WpjCCDL1cmpqANJLXWy5vcflNPr+Jzvkff/hNh0XqO2UqODKuNaTVn8+XtDodBZCuLhV5k2y
lr2P2cA7de1Gl2CSrYKtlKrDMfA36hzx0NdlYhZebjr6MzWar6xeVQh537XfUBpRZlrzVvnHJwi8
3mBoZ8rEKvnTVyeq0leVDzGsV0iIqlRcYETJZKT7Uf4GvLp6ouc7rR7RkWjdKqnjEosoZxvgPA/s
tCraXMit5PGss8Ze630RV7a+DbpWf//znG8Op1mthG4EeUTkAsWip0S8mzkvBjVapAzipDyf2plD
D1XRSjmueXz24oJOV1X2yh/1RcYUlxfHXnb84iiHTtQzjRoKCpZSjKzCMEqbs3MJ338wCj14Ga8Y
gxxGlMuLtuu24ewxRyY/6M/AZ69SEvOOdTlw3IXp9wQn/Otc8OJ9v+CJllWhCUDgoUqTFBsH6w9i
EsWmwFQLbKWHyVgKRG++reVZooHwHwe61K9w+Lr1WpvJIuJibp0eUFAdbKRHFdY0NKXHqmMo4n8x
rzzeXzta5LoyK0sZ7FSUdnXDfqWHdBo4ykic0RoXhTM88BCLF2AK0HR7+KC3Y62XkfiEQwGhFNAk
AgzmJssDaK9fZuQGa2slhhLQge0fkmOyhQQoaFZAcxXylUrWzciujuH5LisYe5tLJVrKDdiruTq2
sW7BkQ1Y7T46D7hMHd39wg9785LsvCqymWabOLvo/vmBfc+Hyo5EHE9B4VjqoH2Tb9jGm/XwqdkL
Afwd1oyAEbDGXgHQ21oCeRWQfd0ajdUJfBaidqCuH6pFDKZurdNFxRWs3Jtsij1zYSLQpfELpTll
72pNGaecp4xgD9o9M887xIk+ioVOcBnlmZLS71XkyLV3SGLYksO4L9hnxT8s8pITRpvndISc2anV
m99u2CXX9oEC5cLw+xv2npxii8YTb9xo2v3t2siyXCkWNQ98hGIVM33fNGpbVUoE9z7l7REi8pWO
6HArzzI65vwSDLXr3eO+YQb20b/FgbjSDuNnDvCFV+MYUilZ++mtbKKp620D4oUk/MJJteLwnYdT
uPgQwVfT7GQ8oUHg0NjHOwoH3ZIHL92Fs8kdMBT8xNKLAsnz5dqZ1tKPiD2OB7RUH1TMzEGT3uYk
T5xQkN+Ceo1l8UxI2Dka7gJJebRY4J5Ie/G5cZmYRsO/kk6rgY32fSeQsSh31gSxtBY2W7Tcnyxq
0ifU6l3HnOzUQzuJDi+gnCfhOUUbbXyAntmW1VsFooy4DRSWTS+U5115BrM0GwkVPZamwyMnYKOV
1usNvnEKLw/JMjI0TL/Q5mJxAGs6uBIffRdOjYFcG+mhfan8w+OwIBICiS3y6jv53EWXYeXd/snv
/kuNWPuOfuUESgBJOpohjZTZMuCGljzWO7aJzT4o7dkDMNRBRPgIqHqdVYyIsrw1tLiy3T1UKFv0
qU0RcEMvSHLrFeGHuqs40qddrtQ0SxZX0/ex+bgsfkrpd4cZoqTNZ/zqEI3rz+M3OCfE/usgDpKN
MHRwSWn9ELCUUotQMtsUuzv4n+KLo43Yheql80hPCKZ21vUlqbMK3SNQtcErGOV1jp9eisFqkJjA
hPu5WA4UMf3Fed0yeqYCShHnn8vDCOoFzm8eZFL8+/QhEa68xp01Y5tUU3OtWf2G7hXjoilKYcrZ
/EpZYY2Lq5N4n8xZH8+X6/mHAvrwXQkPGwN/1EHyRT+G0amePKy0nPkuxvShATURv7dLfzFSuecg
3B7a8Jq+kDL66byl2d9D+Ou4Q6cT56nqOGF/dz3hjAixAGoKMKFDZ0F2gQZS2qyAE8B/5JjJDyXB
iSxd5hGu3wDhZMYlhZA3eoSTy7sw4EFGqrqdt3zAsO75DInZ7xsPsTrZmIeAJuoYr0l2U8e8bdYS
zcb/Uz2XGSkgdpGoEFDqMg4vWR1iBqjP4h2dCiqD97upX2D8WL+Nj9WEQchUfZYjjgnqr29eJrU1
0c/ujtl5swb21xDvySQbacMk6yOd5F4vY9bhU+47RKxnBhl3e7kA3vBfVamXvey0nc895qjcVyLJ
QyLSpd/VAFBoyfly+rwx+P1AJWG7Xvu8zvQHmByyVHxDecrQMHLRdGH8hmfmZseH+uPB15bfMBP1
81Ecv37r3zV4NWgfqJW1NM+n2or1dct1FqjlXy7RQLYhak73LTIHWoI+WfIjGcza+RA+H0EMyRbw
uYBwGZQncD983sYcEHejOaGqBhd2wW7q7gBJ9hnuaDfsI73wCLYQsf4JvkW/hVhYotbXVT3lPf+e
5wh7rhPb5O2gW1sNBXH38ShWXTO6UPUkJNvn2dOM5qKt2intXEe+npOTauROVcwmrk2UyANoqlTD
73wPJEQteMBpHQ2LR1Yj71/bYzyDBWRSox6FRbEpANeyzAGbbLlfx72gllnLTWlRH9F7lOH3EGt/
jJ4LFOS6zFb7+03AvZbPGU/VBBXAcqHwPiXDQusD8mqwncOYGQtGTbhTUzPlL1pqsowht1LgcUdZ
Ex+QV4jQhE6A3A225Oi1XkJDGvXn8T8eDYZI3aD4g3I0PAXLZjEpR6J9CF44DUFBGJoct7hdocL7
buWcZGN0TWxIaPwL4aqptZX8wIkG/cqUsvd22KdJA+wTDE04BGyIA4rv83WrwCJeDlUarbIvHaIX
wHHnVt/F99HFqYKWWU2nqMVNRtDoQKyoAujOfnebg4RY6rgulsrtUqb0ooIv6ju7OryU7LnPsDMv
n896FuVDTuMI8PqGYqWrcZ1QdT8cZp4knk0B/AcdPLMRsUzGjqLGIOE14QDwPiTPA54Lewj9GZyM
lBDE6wqXQ76omXdSs0ye5Of++oD2LyIlOKxdJny/emDCNA2yEmbtOWO328SWeDPom9h2bygSaqwD
9MHuZ93bEsRX4iACwWK8rrSPjaaQ435BP5wVJraWxU+dY4vDlh6XmAQ30TV+J5sJmA+3K3IApbYQ
3PouQbDl6ovmcL/ZO5FnQO4MCjb6FAAuBtY9x6zVsttq4TSXwOY7KKgAgbMWCRjv//5Z2hirMGkb
eO+Z5+oYHT906iHxA05Jzgvy/zhgHIiV08WQy5kNx3LB1Svr/heM0snjH2uCg/FI84D3z7zVMAPU
3rHLhm/cb4XHahkdNg08LvDRfUBQqSx82BfUjjXw5IE8YzA8PO+9slYPY9MbVfUJYQrsx3uBOYRK
+Jm1OLJbOAtEW0zphxl8uDyY3aZjuH9kkMMNq5owRxeGBUyQ6ank1I4/mkTu1yG5fDz0VD6T9zvA
AFhQi1u/RvQjBsqHF/sEj0yWf/nAN72y8TBSxv5VR5PR5a7gTNjYnMwuZnLmy72DWI+quoC2viP6
i/zz87dkwdx73vRvkZber7D8n3mKlEdppdM5VIpEZ9BCmy4knWL4P1BMy9K8GfD9GDfSLLHTaiVa
5dcfEEVoC5qoUdEBnuPQMmiURSB5Xuw0Er8Cmu969KXvFrm2yOwlgAWpsvzzbCb3tJnn5+rkjwxf
40NybDNZWZ29E/7dRFgJgVS1xSi717SrIQXDf1EvNHtT3Hmb7V4UbKwILPNpBO0XkGls6e964mVT
SOkX2D8mSN00d9SUw3cFJWf4PnAvbgW7LEZ1h1qFMeVreyZyNSm7sGTvFGK5jzKDq6jaMIXX0Ekg
n/FSL82l9iTec7ACq3aDt+0d1KqayAMHosZHRbTrD+JT3Go55H3JP1C3J3TbZxAY1gRh+1lb8+MU
rY1cZYjWidvfSl1rkjhmoMOA5MIrC2RlL6xdvWm2CEtj8MNvjdwkKRRLe9h7qtBIHoOWndAlqSBH
sgp1LVshjlH8NYT0+W0JSzMEzLeitJI9TyozqA0cH+Mzi7TLfqKY8F9xegYfYQ2RoaY1+rM6D/zr
cwhmZyEmUhu/rUjARo7rUKjGdRXaiV45w2nHNEWu+toQLjTs9dFsulNv25BMTtAEj3OF60An29bK
L+63LyRw4ASZ0JEwbnpvlL28+hmow2HPp2H5TfQlDTfyHcfN/ED+xBdUpxWl9KLvE03vg+3PuCPq
0DRvRdBvna1uZaEm0Gi3qkmTXsW+FZ97Qe0YgAgG69se3ekukmQC7D2x5GYxz++OFAH+cEcjrNII
QoievK947UifmB1+L2b/ARZAS40hWKdXGel+RReus640rcZORVUt91KgH0ofnRCdnkQg8j8x985J
eoBUCeA+/SZe6oKEwvO9cv1FoRWZIGtJGydbwf3lEtohno/0PECRqeTqBArwO4+5tDTUy6p5quD8
0UcFT/2D0pudF3uO232zIMnInmuit6kVgKCSh1M/uSbGhWHGLAhoPVLfyiOEHfoyH7/C3iXehTAJ
/NGtWj4l57BzRqu+h5Z4m8LActAUPywM07lsvLMTTX6GkzoTsaqU8lylxsiByrGMYAhJQ0YgjPmu
KhnWq39HKVBSeUDeg+9HlYSOXAK6xGIRTu1kno+VpzAgRfEoR0Q2umxetViPpc4Z1Lizu3Kpoh+U
1kjPNbf89/v7c2ST6bAHBZqCZ8746VSVnyaaowB2X9gsatRLksdSdyEow+hZrAu1gVV+rt0xrUx7
7dk60PrD335oGPNiVQDJmKAqEjxXMlaoaHYruTPUO0ArLB7DMe/LcaOGx0S9R9x0Sfv4go7Q2lss
ONEG7U5dADRL1CFzNX55WOYtTBgh8GX0KmHorZ8ghCmU0He5nIpv/VRY+wRkCQIDZrR0JISv6We9
8OzEHSq50EgWpykfjALPgAxuWd6nFSG6U2SZAuamvW3nn0k4vMT2QdtW2SBPfL3YEECkRGOSJNLT
iAAGdW3U3eGn3IoBW2ERhovqWYAh2kKtiIKfNnSKV1Z9ZFrTvdwY9yH+++atY8DiVS8cLafaruf2
cR9cp3BiryEmyhVSR5pfN24md+/0mP81Oo6HgWyZqQ+mzkRxVInyHS1P+wthWxhJQxnbt1yD15kT
8aTTmDEMIcp7QH54YfZSW3FHlwcYXfNH+xib5Ektnldeig1KmNMMUNCp5kmrEpETnOhbqHsrjmkX
pR+XB5ey9uf0TFGXuvLBek+Xc1IX0suW6lMXybobKe9NewVmSWHg97b42Rt3hCoKhdepJw3/g+B0
/EVEXFWnH6cXDqqbiOttJgvCj5bEZDwmLTdgZJU9rRnlnqmfcYONdVM3JHDNDhjKF37MmvVAXqBa
WCxehZ2FL1osYIVhGT0igegIjiH7HwsAo49KXNY11E2iA7p2qM+NO7YTKaTx18FIFUYx+onQwzQ4
B9cNFrx/zlNLa6N52K32piVa337CBi5plOHzeRRMg7K6qS0vfI+EQs1YiCpBEU4b0M8iQa8IBAfw
DZVzDskwbv9yYXOrQKrTPXDdYJsfsZhczrBmbhGEihNRmcV1dg1b59PGUEG2nsNKwhBYcZKj7zks
M/iWCGw/o248KtTc38hE/gpRtvtKyZnk5gNR2NsFFOx5XKLLnAUF5Ks7GTlW1A39YwnNqFZYyq5Y
SVEX8I36pvgi29AzG0+UiX649kQsTpNasOdl6qe7HFzrtg7NPEa0+ddVIwG1Lygd56PV6ZFV7KZ5
fzGuEKvF6b/PdE35x1IntGt88m7dzm8xtm+WQqCb+WT+LQlPKZxBfySvNZqqTQLZp8W5puS9KS5k
NncQfo/r6LuasBzPHnUt+EQNH9ZyeXcfcA1yA+HioshpHaTNyJZwOXzFyH4x+v48P25T1KoOgmnu
LtnpiE+aCrwk+S0f+xrxHzDoUO1qeWjNqLBXTd9jCzvOQexjzUHBL1mUUnZP65DhSX0OKJz3x3Uy
wVSTwtKEP4JeP6HhxcaKkA0SOEfE4rW1CUXaswAeQx1u0SmRl5EPm5Z3iv1ugTU9mrqHPjE4bTZL
+3hfMCVdPjvWF5jvwX/rltgelwKsYnVWfCksp2DdveMBkGXyWp05GsVL4rSkk0ioe7EAj0sJONxQ
EGQ23bjNDKCMT0lljhJoakR41qNLxX1ClaI7fL8zPTFhPaAcZ0rI9gK0slQEU6AzoiQ3V4YwK0je
bwrvTmK5LPPpcEttQenXHodWhb4F77xmu5wgmZsfo4qo/+VtCxPywqDkLDUF+Hdzcd3p09MOYvi+
HDZeGWMpskle1ymb2ZIKliDLP86RfvUbts8uGAVJvFttduY9/f5KdX7xful++HuXPBdsmZJqGxT4
DVPYwlF9l+5/JvSu2SEJ7NHA1lwKlQwBCaxYpk3ALNTg5Lkp6DWqz80ptk8tcEO1vqS+v5+JdVfL
NbdQ7+7vuzAXTgDZmCwRlOENk4eLDlXSos2a+87voo+nsgMILVoqFMfAuohnPnmbZcx90/TM7jZG
gpTyZDxZFVRSsHgx8O8OpbanFOAOEUI4v1TFa0iJCYc3XL5bODfv7bJDMyXGCdyD5ztK/LI9pMxu
RqCxfOCPElIQ22Pst/ZSwHAX4zDKSSlvlKOr9sAbPD1Il6SlV+MrwjpTgt7M/G6tZfTXFllZ2KXn
QQJVv49pF63183by3nvPWhr+4ad+Y4FIm/e+5dg7bxkpQGCH//2hRe45UIXZheGC+eRZjMIAmSZm
lHr04Ch5y2qXXin0JYN4rTKUJP+pEal00u2jXp0jDI/LnC+rdmFBUP4ToIo2x0Xw43VwLnrboXvF
mN43a/NfDBLbeRwxUmKXlsy9r9TCQuzzQDQwnaR8MDIbSouNxWaJpno5d84cf5hVf3ugiC/WfiEK
bdpxI1+x+vp5m+t0JXddxTNd04iPRV20mvoAbdtiMSEOnkHKzOfhBfmzNXGWaAlDQky3BirXXqVH
SjVb7biqj1YipZOJNy0hSIMq+K6WH+6OPtSu+N1Aa0RjoY4xZI/i7kYgBF7XTDrmm9QHIG7NBVsc
7lz/RzyLs2O2qmU2IPLOE5BpY5s0CnlyMkawjqrJWrHSwsrrn1enYT0wPava5ZgJsI/QGBhpvkpS
myjeSjfal0ntXsNmU06n9ug8S3cFdA1/Wphqb+dqTumnH6D/w6e3EAzWs8FLCYNhgsenErQn5KAS
LOmn3cBvFlcandxA5f5JU6k8ZtKT7n3iz6e1L3VyStAURtpkUZ8vviWvPHcXzgtOl76fS+uc/YAD
8ly4NtV+0AY6BDjrKFihQH7DbdJx9/AWhnrjdW7SLmINv8P8hxNaJxDPcpcpRTb4QCAOGU1bGajE
nV7v+GshgjJFTUsQ3IFJaKLkjUS3xH1E7GdvlM3SmxkbHxpRf1WbEzewtul4+7UZQuN+J5Px8VhQ
zQ4Bc2hIGes1kRxrEZAoFMsmrpRL0+4MjQSSVqmQ/sqOHwyS7fCwejXAN8HvGZ7gbkxPjndxr+U/
mU3wUD5nLAdQBqysjXSJbc2E5X327eTU9NHbSArz4O3tPIvBpTQ97Phz1VifxIGUkL8H8KL3QaDD
h7Oo12HksQDdsEKabiUpeegIstjlwXqF4penynsyiF2Wz/sLmxoCVlrR2mGMA7boHx8cDb1qisv/
pWkwdY4kHI5D4fKzyqvfI2EovSrQjgr40QrAJ/eDvu6ZILB4ZHEkMNWzi67cSxRgMKaqOhnynjB0
oqO3y8r3Y+mJEyiGgLcbLJbS0tHntTz5UBBWFOYTHnTDs1K/0tda6WHPZxoWNtIc89vkyINO58nI
mMUUf75Gvhb4lQlKnUGLOaAMg1dDMD9FFuVvqieNzBeVbdVF1y3C8H1yvj7Y0RcxiO2uRWZpQI0e
aGL6rFIuZt+yIGftZljARpstgHmYOsdCza82iycoDdkQFG0pbkRlbieJwTAZr9LUt8WyO+1o8a/9
CSjQEl9WO9H6QRpr5owZoozkFDVpF2/ZWCrTCbgiuztxr4EVjbdyX6zSGEfD52BP8epB0VBwkZoj
iT4oryqWeJAxaZ54lklELPbey56EhHaXVmA2YBoPuzDmop/6hVvIZpsNgtAWrVAyDGqonUy/D8Wf
zw/eLUod/Xuk7A9+pw4qK2f7it7Kl5d42DeJzOomPlHtaLuInrUyzW2SfJ13sL2hrgqmdF3ixHLX
fBznsucnkr7bv25gNryMMWh4vlW73ebbo7ucu13NPsTJSwqKmxFqwnUsPTcXXx+YKDpq2Z+QwCzY
lr57qc0SrbRTlYb8w3b3XuoRTcqSacvlp7enx7JHwDutyEiMpNzRtl/PjRRXepEUg6qkLwPs+rf1
mWqSN30tdQl+jcDJeTSYwetNMrQGmoWkd7wJgRWWAl2Giahaz68QyM/XqzRR7uVKFbDWQWdehKh3
8Kn47yl8bfg/HD22JxVqyqwz5RNDNQCnna5NO99YqbazFtr1jILDGkJiUJtbrAePvUpKgQ6tSErE
rQw20JatM4i9IfjLQe1l1k/7V/bwQqmnONb/3evgSyDt0x22lGdyW20790ra8YrudeOmc+NGcbni
XY4+36nVYd82DMSDyHsyh8GYpl1GMH1NDg9ezArj3TKJZsLlsqLXAbNrh08Wloqwr0ewxoSijIWJ
ZCUu0bhL7LrOrB0wHnzpT09Sc1YKDaHbLxfAmV0AvteVXJHic/rgevl1mNcghv8iGhq7v4BTFsB4
sxYl/lIOEuDcQE+xGJbpAzN4Y70xl0rUC7k1/qKn0/DInvhf25Fpd1N2Bn1Pb5IAZrvUVmUDuWb5
wxj2jZd/ntaVsFxcajeGiLfLp3o2bDv+SkV5T8HVgajdv87K60hcA2TkZfZnNqvXV+DeVXSxxSqI
V1sdg/h3tJf4QhxZet1ZoFY7e+A/bwMxUm0SXo3ATLPmjiT6ooouNu3GmLhqgbySNtcqu9BDmMUf
R6KWeR/hix1L+qkdkHEX+AnE03qU2IsuYYBNo6UQg+TjFRWhtY0CkdGutRtT9ws7HNfNjoM2FiMe
E2c2IwKl7e9NqdiLFUYWzI58YnvTfhf3NnauuIoJzUxDN9sZBQz05wIYQI3Oc5nsYXdi6RVUnnR6
hbP3fzf+xrh0tIA9vr9VZ8qCJAhFV1evj89RyJy6q6W9nPRIHqWBM2F89GV1rdvBGkB1T/sStjDm
rrInzfcjV24Ri+rkfVUpd2aIt6GKLBtaWpbmT2hFcxy4OJDXrb11js0udww1CyZ/BTWWESN97VWs
9nvRvYelwM5QW25zfq/KIVNMmNVPx+Lg0KtmbTVijp350MDLJ8rjjr+6KjuAV7sr/DNghajaPwqa
ybJmN1NjV8Ytp0tKhGXpTB2VWzwMTs0UCxXdg4YSKn3U+BZCD4c91kZo36b9LVZC6loLSSDUAvUo
oo2vdWSCa/vKxxnj4Cz50W+XeBpid4eLu/DBHaW+CdcHq9K3SQQn/wquNgZIKoZnDVAWh7Cj0GAd
py+FZQPGB4ef1gy2gwINHjHyIqc+jI2seeLB/JqzHMZFubl4W31KaP+xg85i+Onowu2dmIY58aBd
viFCmPz+xLhZgLQwli/t+wxllizN/e+LECWK9GOVqy54n1cNoOVUhMiQWpEVueVfv/8V/K8fpkWL
2g8G5eYj12mJdgEGqEXVX+R8eajU8uKnVm85jORm+MRvIS8M4zOVmIJTFCVEXyysuG2y3HshXTcL
bkfyUbWaWn61HUtnd0oloo7V0dOYPeO7vGYH8/O5IWdmFOFtrtv3y6NNmIHziJIuluquwzVBBU/4
89Ti9wCWfaQFelER2AYPCjyuGDNGcJV02uu4xLMHvChe+oqnwN2kPyR3axITJ8oYIApiHaxEhqEv
gY0z1KjWYIOqXHVCkuTUvnj4baH3Txq8f8d/D2H7TvuV5T8kyhHK6AfuM6hW4OuLkygjyqvnc5dQ
uq10OxzbRtgGR945ZcRuAP/0wL4ode2pzGQHWErjENr0WehGiRnHX5d5VFmDN7ziadFgCHmlxLtl
y9l6nawarumwcCCavAozwV2wCmtMOh25j4w3QziUAYp/xYkRUyJ4Wt8zv8qkz3VFmsljToO/AY4r
1PxAb+mlpgi0K6gKP4L7PiSLpT0HkvFCUevlKm5aMMgPrxWc+ky8SuNB2yPTAMmjioC5j9SO8vAO
ZKjBayCfA8y5tPrCW9HkJkUM6+1R8RSRpSuUJg60YNnGHWzqgjrV7kcvic1vwB4y/AFlmGJ/qUhK
I6HR902+5eoXQ4lS6hltXFixZbdwRwkk7u9bGE5tc3xH+rrZqJrBrVqQRuX7drNx3SYGjkcvw9tv
0+jhySqmol8lvZqPoF/oGPX5K1UIdJ09MUaZGJbenOVAYKERgBIBIysyPUatPwfflyYYziEhUZei
kLKWNdlZxhSHaz8UOD8umATEgGjFQEngNdxmUMtiqkTDzUphDXc3ef+YiQJN+yVhPlIpVSWBkI2T
jLWcd98ASr3qTjq2ivWAZ0K357kwJh8ZPv0JhKQiCauT1FBM2l2JmGo//xA0XWuz8VYgw9IDtUZH
MaYBTY+aJE83FuKsrhnwV4OWFVtQpcIEPtSNUlBdSET+Gk0H8nIQ4KmspmTQXQ7Ecjn5enhHKBLa
k+uqgRpAi8SYLqVQ5afEu7Sq6YntueDoOu48JvS192rRJc96S7DbA7djT2gcos8/DWD6HjAuUJFo
FPDViSwmiURD77eqom6+Ok4zGKW7/dbhTboMOBFKfNr84Q/AXm0USG28iA+ybcU3toafH9hFrlFY
9R7AO31Z6aXnFAO/4GMwHieHrZVk7u7DQVYJXFmaOSVjEnNMLwNnwiHosRzMX1/nn7fyH52yBiMy
F74tNcOkkK9Lj851DXii65c9rBy5A6VLrgSiz0IR2ev6gKjjwM+8j6udjmV9I037Cp6wjpkvSdYe
jSkHpmbvpxOyQW8S0F8GKUWjzhWccw6dk3j+ZdWeYGm+yFFGbYJ3gIW6NKNUG6UvLnMYg+oCcrRT
vOvrewh/TgTwNn6rgzBVmP7sSFWstarFteFliEiVyEtUOuyDJIkjcAF83BQ3U79p9typxgKOUgWU
L610F2twEifcfoGq3EUUW/p2MTMgREsqMOkg0UhgeL90+S23IPyafxkp5wky519Vrhwl6itdvkfK
TqPQOKXA8zEzsX4ZPLsmKbMcp9dihKyNeIwHlkuHZ+UtxQqNmT0GGGq6wYrKPlkwnP59ZAaGLZAS
QVXSSDfL3tZO8jyILLZRn99YoDRnn5KXzK66/fLNoZux60vIYsI7koBabpu+Mxol76NegFn5Hc3A
eaR4CAPgN7HyIzvqkGOiFtJWYZFWlav6/PJl9bOYTCLpLaqYsdNfRXErnpAeYVY1NQaQ5LwLNW3Y
XRemAb8hHwqo40Edduy96bAR7XyxkZAv4Ty4btHf8K2xtLFCbAbx4xBy1LBCwss3hzzPDOSWC+D/
wXPL/cneuLRpaC0JHySQ0s4b/2YaCY7MMy85lR8nQlJwckci6Z1rDGStK6hE59lL9hb1bAGnoCTV
eRBZI7ac91/3wtM3syO/r+jr9+Up7U7M9wy5QrKhIfVPS9JkMcjSMRK8gQwSwryKBJhabgc+8fci
RUATPH6doe5bh6Y4Tg7prIcPFMLT9RGCqbzzmqPUFAmKUnyu/eO0pOB1Auyw66o88sLR0J5TJIHL
KdI63/jpi3tr9MaPF4/5WFuRS1oKq1D1vpyiX7zcRnqO9MhbiSfcfT9oibpozEtdrfYbfg4JNeM5
QyYG6u8CECUFht+os+33DqUpNNIQYOF665Jl4vcubGqJi9G7pH3jQ+CXROVTwRCTEEP0JR/dKVf7
j3YZX4Ze+bb8t8tOenJw2V/64uyH+HSqoUL9C5y1Qp+MaLqhfXDpl66BQhFD2IKAFI4XiKaO4F9Z
2Zey9/z8YBPBo4BaUoDYXpnwtYkQxTjIU+TiNslXUgiWG/ozLLM5kzN/3s/hG/zHxGMFIr+FGxMa
Slrra+fX71AZyT2OSukQnon1Y8k3OkxHOAgdKOP0Gclz3PT2FxZfe/C+o85FI+C2ap0NRsTlGEeS
DWdAMRAEKhOTSAbc7/MzPszsAycfc8wbENLTJLrcbUKEoxbhvFHSbffMnJS9BKlgFtaqxwRGnew9
TUxhjdhfyPVxjJlIz242nOSagSnW6N1E9NfQHTiMDjws+lK3QzO4UUpLYCzGp9xzloW3to51Op32
s+hbhj6mu4qoEe5T/FS1dMjkyGaxbBUJQ+P1xEBUmtjdWcPqPxU8OxMLj14D3s3F3U1ndFopYOlo
P2C/kK7oUchF44saQtDN1X7tGL/MjI9rW1L86kamFqds+BCJLyJxC+rDJR3kHmQyUBaGiqUZfEVW
Y6GumaLvAVLZmdz7A2yNTW3rtpRHccGQF60FDFlBdHih1R7d3wwMUznX0U5xbCa+JyGfvc04uJ2T
iJWrdwxZQ8y8Ar+lPKHU4USXltH8h5dEicR69Tg4GKVWeoxsvjftbrwayMLYwOrzQdAOUDVcPY39
n3L4+YZyX1+bE6PptAo1LNXVLgDpnhy3HNrxVQV1s4fzxErA+ghaaTJgds1Rd+1E6I65r12eOkCP
JYf5RFIHEKRDIH7I9TIEfycdCWlRtns6GcHTQgQZillzQn3pKG6jaYRZrR5PNERWoLOx0lG7Fv/3
zsIXWhCIUVwTahZv1Mk09NaAvMxuEw8KJzfnhcwD0gsG+Ngh1YHnRSdlLDVUZ1s5nHQUH54wIPY9
rb6FQS8hJQo1eF+tzYy4vXK4Wq6upZQ+jfgFvEvkcNCy5EaFMmGXyb/tBn3E0K444AEEKCT4paNo
bR7vfjRBogqK+6qd4GdNA64oXgU82iY4BKz8gmQiYy9PrwHrpaCYo9pSUgJ7TU5Rk9+3JhlIycpb
1buEm9JUTzrqtAs64PBFEQMaQ7CvWUzCp/nBT6eEPmuqlh036EjHVJ160AX3wni6M0A07qKosfF2
mKm+8tSWY/vRFdY2EXqO+03hNweCLpnumTXYkuylC34ikdLy2W+h+2HGcmtLl0BOUiAVrwD9fVlE
NbZqv7blE9T9HHZYH/SyKUl8NQBWt1v0oayPZslDIyLxM+SMUCES+n8ypkCUorAF+bPOuEOZ9Seg
yANGJw6Vn/4mHgCd6MFDepzomukEvsDArbWaimtyeS02DTRnEWiHNHSc6cIwxckFYSEVxNIfKiAq
SXSjumukV0j2apHwgi9hZaQUTy3GvvCLiCqI+fDUWIl1FZnnUD9lvyeUR1V/dDarZQLm74b/jYFG
JkUZ+eyQLc3X6pTK/jlptFKOi8pJSlq+kU4tmptHZmqaIzJwjUpgJ/BP+OFsODB8eRDRbXn+61xc
T3jwF/XWzEx6SZ4SaNbC2RdvB/bW9KdTgFjnRDytaHBpdSTe7vLoemKImoRzSXDeoN2+sLRxzSwg
Rouh3Pwbcd8jNzTChxMVD5IHeQYopHiwa2Ml3j3nWEZ8V/Kk8+FZ3xDeZHtzjjwO4oQ+N4OD7k30
IX/qxQZifq0cgkT8xU6ekdqlXVSLGNKr3iXXazfo3Px/XQdj4sEsIvdUqfaoSL93d2NtdPeuoKqa
KVg33JybTQG/HkOa+hXfYZU/PQhAcBJ8uvgzG82XHg8TmaLVXuQDc/QSghKoL8Wn+ZTT/wGoQKsx
CPYqHZpJXb9Xg8Q0snaR3w7WWGUd7ztWFk9PbvqEenFcwENymGnDy0eekjwoViz4z8HT4u5pKacZ
+iBc5jli07kO2iDvnIj9mK5xsGt/3+Q0IuQJzgmk8IPZ6IjdDO50BhEPaRJhKzKXW0yph0eVp8Uz
9ajLv5JBYsrVlCbdPx5ZqIX9gSOn3wNaQgjbWTxi01yKHslfyslxfa/7cNZtRtCJHh/WOzbMfGCu
dqE9YjxHPAbMDr0JW5ZE9hcJaK1wssx5l7+AWIfrf+E/yN7BCgdCoaT0NVQXUtVozereR4joY7WP
0y2x4qTnMA1EEppdCsYNLtW4vj8LfDMizXY7M7z4dO6nb9R2YzWVf2PesdObtmedndLQxgfQOlRH
CaArNpTTEGC3b53c/0Vlm0yoMNW0AOwz9958Y/Xeobwl5yIUVWpxFP9+unqnL/du6FeYV8SaVmNq
0JO41H2wsIdVizviP4Y4c9fU62lMhk9wkczpklrtyA2KUDm36ul/DOJpPtx2w6U3q7GEwLkXiThS
IhT0EuSzwo+bF2vTW4QwSdVOQA6q7hNHKDTP29RwRLqR+v21v6PECMcWcDNkskqxNiDQSUE5BT1Q
7v6cdREzJOT6MguJ6c8V41+rE0TvLCCaIXKJDOYhBLmYM9UtNf/49ae/50/ZaHO0WCyfMEylBshp
34Ql9k9OB9f3+tOxz2V3McwCW4yYZs77fOfyH6ZNSy8aB+rzQrwNDbgEpflaJ+gJZZ6E0UX8BkLB
l2bWDpx/PoftPeTVyE/JEa8ZeG185m1BFrHKwnrrRqKAOtTGRgPFPzswq3OVsSxK6n/HMRy5GEAu
xczxBLCexsaHeaWtMHdDsuKexVl1fWDkQqWvcX5hKkx+NETB0HrGdIEURjMn0Wlq6/6a1eHYMDhQ
NTxaFgZobD7c/ofOBJhqdC1xIqsNCD/gZzN03i6ImKrbL90tQUO/2wOvH4S0sZ/8OGcKosRTbLam
pe8l8nQM+gMZYZJ4IBLAt3sh30hH4YNw6YyHyNAuKiYO1XEBInkkRBlh/nGS4VdEqEjJjFzMMqlj
HmwpG6acPDz2DRTQZNySri6qLJhJPd4GK1rvZqaHOW8AIIl22zNgTX+8XX5j//Y1EGHs3ICRFjI/
rVVSXRzpNl73FJhAMOlQBjRDnpC7Ksl55zx6DbV/759nyU1s2WIqHJ++M/vTGzENpoU3HDsUOZT/
virmpjOmD73xG/+NimPKUSfh6KsgViR+Y9k5zglqs/WBJs+fE8UchEM/B1PwwIhATYsjuBM57iSQ
Yn6g8WnwRnWUjTG826N1t0eC0qm3oWoOEQlEVqV2szUz/9QUz5jMzcFDmoINa2Iw8jPp1V0ubUOQ
z5AHAdalIUoZSxg4g9qqWbzhQLvgx/zkGVvc9xVUvyXPa8PRRaxC3qd7ecgMvdpoHuyLVN6fZ1+9
JAvmfpmVOmDG4UQufN7wbDqL8dN28JQ5JQ9Dh/XCtiVOVQS4Qn1gSTblHcKsqZXja9kG3JmGx10Y
Kam0ywwA1SWeErruLJcUkCPVOSrPp7/hrrPPRwgjj9Lvk6z7tJAFW2W9+9KTCVF6kdhjh2YCfZr+
QF6s6xqflS9Xiyq2TFKPl//chTVnUwdG3xGK4jWra9HrFA3kK9Fpk6WlmMe+gOwwZ72pf/Z9W2x7
I9DG3Shj6+KgRkj+1HAzmdVn4Pe5sJwwHpEvv+5Id/VSG78h4w6flyBWFAoEpTTLBCG7mRTAHANO
K+Za365x34WWmExeaMe/8yljZ42qJJJ73HwUbwvFPv2WCnXarEsqP5zKzgLuuEaCKuD60LzjQHLo
thNKIO1zOmKg5/LFwxUiEu5G+kI+SmEL9NhhzyLwL7uLyQ9jQCDPEvytHvE6FJtkYB5bV8SmYIyq
YuNGXf8a2GRwJpX2Nw3vMgXwR6qNwCTqY41dt/GayEQwGYV8GwuarXQCf8gCfTYKIgRn5a7hkPSE
8ezeBS43En7o3XhC80ALezk8IK8QrQ9C/bzJ+jhqbK1CfHdzFSjYaFJrkJM0cGLu4ZeSRjbF1jUD
0p8uGy/xEmQi1Q3d0AmORgw+677B13tQtJdi+Pu+9ZaFfgG0jqowno+1wmPKmG3SMqGL59Ni8Ylu
3pHqQtLMiDp91iP5qkHsDpO6XF0BhN7GpVNyO4ryprnQVEa5GCUhxIlcw1oZEjWfIgLmIwBipeuq
awVM3mb0PRyc0cSbVfu7pSvIQoBIblxAqagSApVE1DoZXwWqibGyos5FqbS1R3NGBvNPQBmRIBDy
K4isWlVCycdQMY+xnlOW6DWwAd3q2mzPRWkJebKIz12/VtbFh6kIiP8v++l29JMsjkC6/StKZG/n
sRskz29WOZatA33FBVsd3vY9wHdFS1AUw+UUwVP5Q55HG7iB9yWM6bm/+47cdQJUWos9q86aQCE7
RN6pjBe291YggJcWCuNy1eKWS7AWQYP0761FPOr5kMuNYixERkxm3GlSUtwVqlkYwAfam2iHWIlG
/iq6qU1WH3tudxe3Y0VOM0zpci3jgmkIILZnamj0EgMWCT5U9cMYqOqPz18UkQ9TsTRvfUQK81ev
X+mA8YfBxysonVlK46KymnYX099/oGXAIV5SlZx4ku6YH6sCUB+cxbs1PS7mLnYBUiAlk9/kMkYp
6jATP+2pc/UXQC71BC2PSgRKBsGRYHFZNuUTz0Qt7qBEtFA10UaOwKFzMZJuBi/dt7K7RznO/erp
z88pUTYHAsrNsMNKp00m58d+CP5AxE9PfwPGsKFIGDeEwMSaCwZSFjQ6i5kZZDcKX1LGW+z+44cw
URzQOi93hko0JFqtbY209ifRQ8wpgUZURLV1knYp+JEm3oxKSQAm6koq3xXWVsLmpNOU2rOMmF23
4TxAHbTXSEdRMYAVF8HpXKH68ceRj373F102L3zGWRu1Ti9+y/KVKDfMHBxwzjxBU6kaDAiylV4F
4QiuFCKRHLwV+ieEnodaWUZkSvObztz7eXXaKtFvEG7mYxrX8RLs1bQN936pqEIgeCXyb7ni9tJt
ZauxYFsKnpTjLLYSqOnt6Jcof2eg+qdls2WeCRusbqw3TYFsEI87hx0vspn22LlRPMuSmZNtY/Ki
UodrnAM7ITEkMXHcmem1h6WLyn72Lw8kf72C6EF++waCWwiQzU2yjbdAqmc0KWrYUmuxCeDFOIQQ
3AWwFTKQENNTBXLhPf51jQMQ4eCgLmma8xjJXvvy1AJGXfUSHsngoHItM8aktQDPmt76Z3lSbS2O
P0a/EVWv8GnlEr5ptyAV/M7X80byjEP+DEkzzSgAoWfLjVdZjWLkpZ7w7VL5+BJSeiYVK9z2x/EA
/M5qwSOhq1pMUwAzWbQDx9P70AAO8pVzuPsBzM8VeJ86a066yWfageDF+1FgOFxgERoR76GoPqkH
eofRP8aCov0wbIOCHLZKzNoDwckCp4QQ3YimlOfesm9FryOaBLRJ0bvE6XEEf6kIhixrxuPCM/0y
M4bfpE5M6cPI+8zI8oUrZUpoJaGhnYYkAE8IBNhk49wiKdv4wsYfKCbEBE3MrBq6bC5hn3y230+R
mZrM4dBECLMKiLGcNI6QHiEMyCDiLy1QSWf2S40N93jBcnC/uXUnU5YXY9zknZW34t+UznZVt8PE
DTjdDJJz//+q4xkolqYSzQU9cTfQ/gigKoVxUWHwl4zsGu6DY++ZaDvtrGupT766uH+tkj1Bu8Mg
iLbu1Xj4LaLPMNUgUDG2hH8Z3ceOMh+C4+aXEadqwY0e9PeXxvwsyllwtAIFqhF0lixNcq7P+Ygi
92pvu2fj4DmI9262ZHu3Tc3yxfEgpL2PyITe7azNr12RRj4fT3bJlpGX6rglm03igBKh6Yr29451
mcPXElLTne2NCnne4HFdik37xhLNrE+vDcWbhtfmsZJSUtZKN/tLUP7FffKKs9m8CmLhwhAQ7dEW
EUa/g8RdDxZjEIOy56mTSPmjCh+djd6keP5E2Ov2VjvHQLvNOSh8NntgC1SEguZFCSb6HQ916HMG
Cbo1ZFTw125f9ePTsIP2wvzPDyFao/qnYkS3anTJIFR1nOyxqhXWFRSw5bt8Z+9eBXbxYI9NiM0g
bw7Bc4xAsvwiLG/HklU4HGakgOJ9HVhR0V79zOzh5H4HsZaBbYGtxmkRJEYkQprKZY1N0ASvO4GK
dDStGSzEVqisajih921JTBgsmoNHDS/YMCgcKCUFlbpma5rSakXaAFLdVLG3k8T4choASzsmUbnQ
eutGAiL2Lbo0PBNqAeGz6nU79PnOOgDmhFX8Z0RTfBpcBcacKBlrkf8hMiuQll6eBOwGJZJ5PGFD
QcgCDqtH8kgFTu/fZcmW9XdLgsChgY3D9UHcSA8NE0KAsdO7MDPQBL7rHDUGI9jIF+EnSuZ4u8px
zqnoqtufZwBvHTZxo1Jr6CrJBD5DUbWhgp+2vAINb2JcJauKsqmB+yNFJcF8faugnFDwMqy8nCdz
gnixNI7qVf9CaoBIafmLE4cvUAK/dt4m3oGXUl+MWFSU4KwazO/peKdvWnwbKSFiNM/2a8wXvPLa
6HOQev7qIvjoNeGp7dLMQt947c4sGUgu9cMFetGNRpwIOJadXJtCalEyQyeRi9UGrFgvH20PRZd/
nuxvLdabBhRXayKm8P3AD/0ZlliNC8ga8OnKkazpDZnkbClq5oKq4RAMjbIdEkD/PGaf4aMv7/sE
AIsYoPvvT3VndWdLUXD+yaRFqr6bRzqSNGuB1Pkf/1uxMegG6rwiTbifj/kIDI2iAWQO4P2uKylv
yiSdYkFAh/5cl7D/jY0x8T+JK7+69NoqEzqmGlQf1OKZEaKZkTzGSvKydnjPej4+l1FQq2sMGx5A
8cZPaEDiVHzlUB3KxYFiyPpnwgF4TdR3bwHQuiIeE9JReQR9jfG9ElLZD12w/AOEIagANFolBDS+
LB/MjcU98+MRMGS6E8KQ+JRinOpF4xr067bL8TN2Ws3DNN8aIdRZ7sJlbTBUPWW3qifuitKw1fHD
s64ixq2VN2x8DlZYRVffMeB1R45SidLtbJ6txSIcD5/hfbSy6QoPqf0IfvzZUrr/DXfBPct8/tHC
Xlpkiz9sYkPfXnwlR3myAcvdJs+4iM4HXHQvyYnib7WIb2nY21RuQvRx6wBQkbNbCqWZPULY/ZnN
4SMN4gwqXJoscRAO+Q/ZGxz4js9183gn+3T+6bmdGzAcNAUL48CibcFy59Xhb0m1EQIIoVeH/TX2
op3dEM2+NCLGeeZ6FwgvbQATS0PhUXgvUrwQwnud6fFQs7MVEbd+QIQQFi7ji30+CPszP/YyLAH9
mDw7Z+BxLSwXDAV1rpz/e14FnlxKdyQEZQ96jgQ1+IUK0UFh3OQ+f09azMRHYO5n3asaWOK+zNGC
FqJBturgcVlqO5ZwNO1tUhZthjthMbAgaw9uukfU4lu6ilBlWoARK5NvH0BqT+yx85DTedPPZw+d
Q1chILgDjkngqSXOLjdsNDp0t43iALF7UZovMWM/i3jwRe3P6k+6swNy82mkbuJgfHbw9fhEOa0q
eQDblOFwcpdRBf6PvDCofdYIYDe+L2dLC7uubm6lnqnIDFsx71O21U2r5sOe1xv+U1rsnqjFhGqI
DZDwYqgaiTa+HIKg5CcXlQ26BmGgaoPaj4b4ctsLtTBg2KqnDbzCGKGYGMeluclfAbzV1M2KxVin
WBYAVQcleoMo8iiYq7yE2FajrtzXHyzbSYIWSO3Wp5pZp5pJ6HXBfJSXhZlXPd8dohT2SQjiCulc
wAn8u/MFAC9HpdUatRo7evMOBbz+gNDnDc25wVVQZsRLaGWnJI/eCs0FPIkq3gaBQTN7o2PyWepA
034iDj1QW4OXY+aNd/N4QgTqfKvI3tFeBEyz96lhkkQ0WOGPS9YVGDed7yYL1THYq5MylWZchBxK
QvHoufVTi96VCjXtr86VOW1sZFGEkBqtpaWEgHzPDCS7tWUuV8vEqMHV6NjmiDDxXQUG/vMPP3s+
1kVcw+3lzmjLnZdAX0hYWZTrqQ8V16k5U7hl1nCn8x1Hcfe70o+LCrtsOkdOiQhzcmdakwPL4Gij
9d5Al6TEwAVvabIf9wTKNlrZ4lrxUGW1AtWOWN5EEvItzkYiWxUCCVRJiNbp9Q1S1ZfjYnfbIZXY
utQNjmFV9/R0a8azSKVxlM+LGSacvtuMLVgd7kBSQJKQVfjI9AhOkFAk0iEax6PLdM/msIGeHNbp
wRdpNRp6DWlmGfVSq6Ziii5RHMzu/MYdljjssLi2YjV4d/Qeumm4FxRssWx7DXaXD2DkWiwwUowc
xaJK0yu4/Y6jZ9GqEi6ldP939FzK7tjb4YSLA1FlrMzzIWTyFBp+NBbWGGlHZk2dz9RNwyHX993o
xR0jEdPOE8pgGmP/XuQGAZ6z6GC1CuPBiY+KRdtsyMBgzW8teEMWgLs3rSSRlAy/ZdYxMg0XrZ4a
nHbtopAkZ877SDYJafXmZpFN352r3qqWM22142zsV2HihzSEnfgDa9yM3N42IXjmhAECEnabY8i0
KNzKcBX2o8JGXUu9cOzpYF81creHbeQqGHsv5q8lJrhsVFaqp2voofOuNExzsUU4mzC6Yw/2FEs1
LKLBQkEqUXZNSCHGK1o1x0Gd2DdvxQHdlOeS4KmkjlRzs5EhPhGmKmL+e1NKCVj7ObZmqPIv3jUg
Bxw0YGUP4Iln2YdwTDgA56xI/C8Fk2k3n0WMwExjGWxKlsDMTYyjJryQrdZ3/vKSk7xxQMZrmtMV
Xd5rax1vnqJTqWTMJ6OvcHum2OU1GRa43481NlpFRI/qyXGoewVTuOsYKR6QXtFC3cwaZH/lui7S
trLkTzk3pzHMQsKQ8zWN0nMQL4cmyen38Mkft4NNQIhBNX4Khn6A5cnXOxWnRZ/j0AUvpuTMVwjJ
kFM7UMKJ6kTHWwhAtk9RQbKsCaFbTa/TRQmLrA2DthRbSczYWNTH8UVfkFkk4lKst3/KP5+Xrr7/
C4iusoDYgBm9rA+QGx9oHMb6DT0TA86lQ9nNS5Q6zvw4IpCRL9ik7kBTat1DHTGAfO8+g/I25YbW
IJOnbQF2IMgycioMy/2nOBpeIch2EnNnoz6JYkplFJyB1iRWCUWeZSU1wTdOfAEk0Q3zQSAwWlkC
u7LKOsRnp/hkZ5lqy0NZwqsK+DQx8d3gS9w6oPu52lDVnbLCVAz+Fv+LT/OpUiUyJu0uN5/iAj+a
KgtqpaEud6kQJI5qbXS8Xm7xoMMAzkolu8dsAI4GdXO7OwrdRwGAvfp1iUq2PmfvkfHHalmgvH9+
fT936j075gdcrXjnyOoQhNgnrIPJgcUs9tI0wO+5CQkbkummDwj4IWRhkdvzmk2HmZmTP30sFsbB
SgrqYzxntzcjRVUeSoNatMQwhJOmAZmxI8f+atuilmfTDitutf0hhLzkexiu9MSKVvzRwvdUSFVR
GYtMKnCZtBPIE+QJNJD1SfHoblkEZmo8nDK5bdIFtoJ+qUGJId4g4wztIw+XR4FaeoqGs9HTLmfp
+YY9CYgMpbrsBI4lbKD55qaUQpB+UA2TJ6qhfopTWkeNp8ExGkE1SLTuveov3UIBxkQ0MTwaf5PB
jKNvnzLv7AtEj2Ngc71Rz6fYs9zfFUlC/79Kkeh7S1rw7vSBO9q10Y42ER5QwzR+P6yrxiycfjpV
/xi/EzpdQG7e6pWZXrsfOZkmUvlchtaNHyIpbU0kTvvIYq+7vZr2H0BTwOAl1HBd0JYASJcruEzo
yLsYUcsqVw88m5+AKLrS2QBFDflalRl/Xl6h4g6M8nLL51CqSLYF8qwygHUgBC8BlULY8lu6qAng
meA4XIS8bkHvPbyvbXdpBOzDDWPYapz5YPf+UK0B1TM+CYnRolY7JpLm+R4iOV02zugF8WdiZgEm
Xk8qL2GRGfHmJ3vOeRAxFFU/wRHIEDdR6SvgAyNn0G2o0Dd3YP9cFB/laCy3mFT8ToMidI4juhCi
07yOdXFL16iO3Dgp5o5L9vnjXSWAdTgRMAEC3S9U8vBH4om2BPIF1wmE/f+k6e2stNU413TVXjxz
yVSJrMBBDNRexiB4Fg2CfwdMrKROA8PUm984MCvddbEBqWJWADJn7D0hNIlD7q9vvsvl7xOaNM4l
dttE5lqykU3KjR18jNaMqy9b/wtgiH5Ld+6sC4WYhd9pVNJUP/6OdBC7PpI/4Y1xFP9G33q//4u4
dfvTbXS1TUi9/ZsBEBssO5rzqI52X+I4x46zarvsqnQWaVItmT09xgQc2WP8U1vOsgoxMQKyT8t/
HyyvNX3ZA5teHS75k/lfHsM4FMVJIoILadxANdZhPhupPXOgmJJpaMeMQSYNXPEv8/OkTckk9fl6
UL2Feg6MFJF9F4Fk+tXSZDo1dsFpLyYs0YKPBInMXX4e8oqA/XsmLn2wNeVgHGujCbcbM42kh+ei
rxGiMVWeGMcSENxGlBYU3OycWCeHbvtrXrnd/Rt+vWWaRBAD22HmWq7Cx4K6nhXGtZcoTff5Loo0
3yWJSrZQS9nmDACr4xqqdSNFJJfvfAm5PazGW75TELREr7Za0Lp9oxa+QXcZ70stDuTB1K4XEj8C
ruMhITXI/zd4ZDMNO0s62Kkue8SVvU7cRZKkuDH/9TcNhrZMiJVIeG77eOutqL5a/oh7cQxAodx0
Q3Plq+n6uS9NrbyI0/tHA5wVad0CbBAeK47w5z3E6rgD1OswPubpmMTWk+R/3qEwgnd5zH7OtQG+
aBZkGUw0R21u5JVZucxvMXg/+g8pJQKApZDehydxDPYZ5z4IctgIkd6WffXzkQm2rKKEida++IcW
WMt63MYTufiQJQPv9XiA1jpoccBbES2MYUVpfd3r9oo1//kdmSI2q84E9R+jJg4AWp1Bq3NMBKsg
DfsYWDp5D+ObPPaSYCOV8hjgaJP58TT9q4i9YSHYAAaRyU6jCBquIyGiQw81VQh+eDD2XCsbGLSo
3Q6cpsa92Py8uac+EYcbuiCmz50BM3hSQoXedtmtNe66GL/OUR+8wwaZHbal4/jZCrBNXo+l67gC
FqGHAHh2J2/NYvOBEXyK4UALOBsEKt47WKcsfg1abUj+vB9oLHIxlRJ7/MrTdwV7hHh6sXcZxnw4
OgvTG69LYqTDL5LrCCN7tZrWtANMoo94YGMZYXmqqZMrpFddVdHN9QdkKms35yLThcwBQ0U9mUok
yFhJXoRudCbYUvGMfw4gTmCSXS5zVC5ULRKa7iOKW97M9TvhwXIL9jmNnPrrpcxxsnrkMDCtAmEh
PnkxTfATa+qojyDwV0HFaBEH9h+YROoPqn4mlv8hhZ3YC13mjItKnzWsCf66inv6qkKRBr6CoGrn
YpZNMqdbiQAYAsuTr9G+CFinr0NpspM+WM3Xc/Jq26GpgyJLc9cX3IGIKh05bSyz2Ih1KiHhhLym
BJsJOniUPxLPBPiHNm80jPMBZ1bTBTFrRx8gAVca3IhFgRmBgDpqPPioZ2MquciPMmgqAzv4SVGZ
lw2ahSNEVpgfYN9cMd0lfhFbeNFuRfnZjseCSHYe0RogAHAlupw2qSmcKqv5r0npv5OOiDTVTsqM
34Ypp8CU0y/2qFQR9XhdBz0sxlsbSbnXeamPpT9hs25mHiY42zz1sebk0n66pCxhVxKgP2i2nabg
7+FQyS/gJBSX1XP83IXKxdoo2tLYu3fs2ptKk23q5xCRpiLndYwTVFnzL2ZLDGBKnyGn78n1pALR
328S3Qg6mjbj5A6RPTGPN6tFdf0YgTPMN/6UnfV85fVU0PrTeslLDfqnTgn7tsZoAL128S9/p294
/XKtH2FgT5IiABKQq78ht17NRfbA6isB4m2sVe4gWrJpNP9zhsB7mWCPJ2W3lidlKxAFDsKPi/N5
bDaHfyPfOhYi2kTz61SIR40cgw1q8YoR2CC9oJyTVNoazcGpGXD78tj/wAJABp7keC+PQgMU6UzV
/9jf2qk/6XDp/JjScFxox7jaYUr9k4EzBaVMuWEKy8yO9KpfZ94nV1ytRyA3QxR+5r9RmbghHHW6
8hlg4fF96nE2d35HsEqm4JCwnQ3iAfGlmHnOIHSuIqlCMpF4zJYEJZpucXO0xl7fWQFqmAIq/O9b
gL4p6J8BDttz1H+mfgv8dWwiZMs4iqD0wDlOdZgEPIi44UX1LVRhX3CAowIcaiMWsYWUzMyeK2Ew
X4I0vjd71SauJXj/YBO4PNdKCTH36GVNO2lUwSD2olEpS/3iLpAGUwnK3+EoRsBw9f2azPLjRQwA
K1BEElXxpKR4yeZXSltt3We6rAkLOf1SvdfzJfdvGp2Rha51wgduIZh7DbZtxad2BDF73A4E6vIy
n206Ia6iADhjaPm7NyaiHDy+cFYaCgAwn7+Yjl1e0naa2HAdo4teDp1IQZUBlA2VNqt+RxYdnUSy
x84+wTh3EDbfq2T6n16GPvZJgXBHAuuAGKncxAORhMaFODIDQgLaxt8qo7soP/J/oENqfwI58FVH
cOMsPPHmE7+c7CqqDa3SsXyRvvncE/iulGuEqbhlmoLw5Tch1xmynrOmo9xZX5D17VlMjYK/IZ36
3bGWuu1RXr2W6xVQ9BkPGWCN2+XAxmFWxihSUOSNcjPQrzlHb0hCJiIF5+hC15eM16F1zujV6tXL
qN70dDqxyYMeKf94yoxk3OmWkS6zirGjbCyNw6uQ1qdWbpn/fPSW6ZQ5WjV385uaHj0fU5Tr8kaC
psdSbps+tHs+pAhIfQ/JlBcG9MrzWJD0Mjg2cbrDVDJAIgPSuCnIpCFPYvyx6ug6fk0euoe30iMp
fFVgXzlqfRf6ydGbSqU0G9QTHfls8/+F4/wqDFrrDalfgjaD4HPdCjuutFiAJfLvoGY0XRAbSYZg
3bn0ExQT6oawM0tvL3S5ZUCPKLMwXhOq/6llfqfUt8qvywsQU+ZWZae/LFbPtuvjdh3C33QzPvjS
Nx6VjkuriAsCxbEJik7C0Wza1heJrEJt89tk2kjocdOTrSa5VMKM2STvYukOvwItOrvbbzfVV2pf
eOF9YnCJCSX4K3UFkqSf4Mr8XSTmjYzquOk26DcmV3pCAqACA0VSq+RTXbcHMrfe2pPgKX8LLz8R
CPSmkpgSB2PiRB5nxsLak/+YS4epGuZ86VUFRQLoAAX8OZUqp/tGG0lyKMdXDVIyQSwJG/oD5duz
/pKxQ4dp7jSv4cxOdu7yNsKzHa7EHzdX5/wNu2KiGgqi5oGCc79o7GLShyCRrfTREzK25e7n9Kue
0G4CzV7CX6F/YMFS77FFJLqplZDcTkFE5nfWJMcBnVUhMwVbHr9FL62jMaFs88d2LLuFOfCYlG4u
zWHRriREa3ZaKDZAQbY0NbOJhNqgKSXq6Y5FDFGiKbua6nrdg61e9eDX+E80zSljea/pCPd/ehoO
r0JdcrvguSOG98nu5mAUqVbbdlp2YpuUFPgi1/b9KVUhPKOajEwJHC4d2LD9/YhALDahyhVksy6z
tIwjn42QasbWgjJ77u1iDiwkeLQmaAZo5fqK67S6KJrzN+cqZeX45JT3AORqoGWR2BzSihHLSD58
0CPIyVVu7Ed+YQ5nAk9CLNqyR7UPOg4T6MGoL3qK8X4TTLlyKKQoA/N7WFTa11ikjZ2OrNY713ES
8iM/Qt+6yW3uhufCtOBV0V/vD0VVTGC6lLNndGYbdbiJyzBZxLQK3E6GzDWaCeY6SvZAecQHSa+y
OEBgqekGPc59tbTDG/BUo64GTXMNSYwu9Vek/uNho1RHLAxTByVVfLbqc+egOqEdbRAvmSdJU2FF
jPS1RDpDZ5jHxLbteH9T0baPUgMEWBZLSQEx2s07HvMoJ4bhG5CFt1Mk+qhgpskr2MQYLLlpAe2E
PD3IZYnFMnwloMlC1I+oJH47J6KE3jlSusRRxstHgSPjTPiOYX/KfE242kFrcfLk+2Yh4+tWVXtQ
J7uGxzQQ4cPTZP/2a2eC2fs0vtqm0KkqLdcmKMD5vaMHTrHqEajFlHf6TjYl4vHiJVIHmnSDaQpn
uB/V8wNg+Vr6JpAha52jLmOa+s+9rbxwXFRzMRnLnPYqB+NIan5aP65sLqyRbTbbREn/NsWGfKue
K8CudBIxiUIMKT8xDFGjH/wVPNUgE7MxoXo/ToyZYc1sdvCYsDMvbIkr2OKGSM2gnRpeD/jr5eey
clZeLw5C6wiiqyyEAjaTsqKw+QOWYL9kj1JJnJ8fv5ZcAQUJcW2WZOx3EGGe8fVJWuRhZx/8NsjN
8OtUps1ocGVrY0jE2VbB1OPZ9H+kK+vogtJnMYc0K6S2L2HXpz6PwS8jrh3xO+KeTrPT2hDT54tb
NpwBfARmtqJTPkQBcDffpCCHmqHGyEhPD2gdi/eI8e+EpHUXV8OsGr4PlonaqXHa4xlNBuLnZ+DD
WuyBDo4cmMMNWO2n227jzdLfZPjNJhfn0LALHFwNYN3RPOznW7pY1dDPThVg2CHkwZcyH98XuR6R
YJUUyDj4AVLS887sHJsxbl87K8mmFrERIJeZBePkK84Tgoqzupj7J4LwzyhOcEubPyVrZ3E5bd+g
DVH9kawh5Ml9qFRoBE401krLN80Cr09stjjaNH+V8203ft2siqg832HeDMQgI5B1Jmjx17Z/UQVB
gBn7SmraGSGgglV6XkScG8YqXqHKAh4ycPCQPBz+JAivCJJlzWDMc+uD92tTfSSoswv5j0jfFngF
fP+FHkqBejSD1MTLAMKgSNduYc/T0w0YvJyURBSEsJmtHECYYOh4g4XrxXqeSCjhJI6FAxTCpcGm
4sN8YNE2vv/iUK6jSdKYCeZ5gs6dcWq0BMQKfW2VhLFZc8dC8KOd41Jx4LKSKkyrN3pLZbU03W3m
ufAzYwoLDklXBX17pXnthUHdZan01RpdDZApQYDlBX1CvYZM8YjxTOWhM5O3N5IE1t6LrAL2JEba
FjS5MFx5SHuPUIHpBrQfTfz50HdwOM9RipNm4d2mxQWrw5mPBwWqn5oUpZKTuUf+yI9cF5OUPIhN
g+BixNhYu6U/x+eDgvyncJ5BJiMcaBhA9DR/rFd9SElh3oVQQrUnxclvY/QPTmhyrbYVbFr5BU+L
QcO4KXy4u0TcBK0QGVGfULKsagMNcljqaxKxGEP4WqcUlLDfqRqZb9tQluEMUUqzTK0lYqpHh2fh
Q7/w5rhF3522tkqgYiZ/c/VAKmlzjSDZd5DmMvrNs81sB4nKpQWowA2Rh2d+PxJg3DGNq4y/YsQr
FCLs5YasRPNBvQ8rztp0m7tcE8D6nuwKg3pSFTW1aIn6EF1JBYyGExQkE3XG97HLsxEOQQisQJi7
V/6tX8c9SwkjdshDwkj36mN3zIP2glzyrNM+xVkBhP+lGP0Q+5XFyDwGIkm+tEM//IVKZ23CBvxZ
2BdFAFvu7m2UDYRvTPMRPrvXQ33OyA1mWDYR6qGC1L/Q3/0RAaTMpKFHIjwHj/FwM18BeirA8sBM
Pe5QDTbvV4JYXQ4YR97HsLvBoR2/UgOynW5b1Zgq8+xX93bqgD5V6IZiKGRoN546CKDO0MkhYOiN
PMPLeIlSRgnlyM+pLx0J+Odtvc1PUZCUgrGO9mKYHTzT9AjtxOftc443UKOnFA6g7VtQX3pcidP8
4Yfz62fWehT8vJRA4r3/4Ty+XRujrcuMHfcFQ7sBdOMKsyk/uZarqiw+JZ2rgxkGsp54Y32Y+2gm
A82uzQvt8rD7042EePDoIiagHS4OJJgl5o0+VWKICj6jwTtIsEJi+yY4kTUKek5OrOyx/CYoeJsX
JzyFcQ0s1xWVqUpw580B+pWx1RzRAeJP6eM2Fgd50zmaXd7yPPXoTVZAwSWLXsRSvc+qtyuhpKPl
+PPfxlVSNAH1wB/WQIyaYm7xQUnzbehD3u5kIIt8OahdM0j4LDeGplHfrc6f4fopRkYKDZAqPbyW
VKW5pA3/mSVN3X+0sJQHsfZVrqfP/SwfWTNXNi4WADsXJbm5EcrERgoGFsUhA1XepFnH9vvK9Vkj
dug9xx0dULg7UTK4N71fBqkABGt0DwOfJ9xlinN4BaLHdx9txhXySrMtnC5NZn9s+9/JtUUeCNG3
z5QzhX2iMdcN1yIxAqXbaR7PN9NJYmyDJpYx26uiVrclzXnKVg+C6lrKcySHb5awCC94qmVXyA+m
gICSnNEDOCZSE2ovYPmUsL/12BqdJA9Jqah/le32cfMDMcge92Zq1mXn/MgvU6rWgCAs16wWx2MN
aMpF68Xvn88/igzzLcZSf0Z/ocuXiS631/6Q9LniaYHm9u1Uu75BRbkz6fPrS3kbS8rC3AgTelOF
RHuW32Yj0z85E5btZLC6obe7Enuh0NZ491uIc0JgNMKNtA4BoBejgSj9o8oCWUa3evvaf9u3/loq
busRfw67/2DkqXM5+K3JAXTqCyEREnFm0XxKqdrHkvXlPF+a0s2oHSZhfAHuOpjyTX4PQiNnniJz
bOdQYGRCVDADOYdrltMSmq2uY2WGsTOjfRSUeK0ZD9NmsRQL7TPyXuO/8v92j+Alv9nhcdduW7ad
lVBL40OS3XYmI/sZC1SQE0KGGU57PnlJqjadbCcLpEHHUxsFREtfJ186pjrUmlP0Lm7tlEW4S2LW
406XplZAmLF7pbl7kHIwu5PRaZtrbfXjDMQem80ZafuyQNoHJDRKfDUiUC5sxgzE4sZ3jcNexZqq
9sVJRuibM98glqoNz6S1qXcA59wuGLAb4qLi6aT/Dx+G5srQj12J4ir8duLUDxMjM9wCVRzq+nmp
5sEduNgXUgw3JjV7Ohvnt5p5SRnhW1V0F7L9+KnAwYcPiJdwnNXwpkGbPiHTcshTNmftDDQomXP9
T/7aEG5owm2hNx05aEn+x1fxXbhmA+Iqe3dzI7S+L+EIn2yhJkNmiar/Rimwg68sphgHDt9xHBh6
Y2Nla8RL7vzbaWjazunYCx8Htz3IsBKziPyQIhwDShFg2MZk+a/d5YGTeb4zp/izXjUAwXp312Xm
20xFkhUmZTWPikTa+4dtKXjHyiSgf/1jPegTqaDLivAWPh3lzbP2SXNbjJeAIULk5/at30pFA/WZ
sdrS2qYLWAXE55ArZmKy8cL6SFimOMiZts8lQgIAu+esG9VHDr45Ojav7JFQ6pDTsCU1QjyhB8dA
C8FLL1XZiQ1JR9PknnOf0WWeRh2hwClBUywkzgubNVQC3XE4GYsZs/d33vQcorgX/lUH4KKoN2as
Ko70WKPA0gYziKSPXDHj/1IRDFjcAJOUHD3Q9dUK6Ka8xPOFXRnMDyP8iL0jiFg+9dSb6YiCL4lp
7YYemYUgXB7Erzp9dfcyvbHRNO6DZOt1WFx8uDRFBScfLmQBNYT4L8BhbFfg912EpYKMMakTb5ZM
JBRrx4zYUfNkJOIW0NHXE1A3DAsRZv5D/oLdcgcq+rCyC9p/WfV/11YzId0J2/i7u9rcFhRKRgFI
l5N5jmc5vItgfchFhGsVohBctEDiFh1Oh8GRjqok2gFdO141jPqadSa8Os0MYWgBstcOdhK2+Plq
pqLfmFwvXg5ZZrK5VTRYa3pRfgWzX306AqN/aBYt7JxQrnGD8XyDM8ImcObSAE/tBZ273fH2UZK+
al7nO1mIWnHS1xigmv+JwKWbWh1l/t+RXm+0bL7HNqJYY0eUizYtnqzBK1PAtKl/e6QeTZ+m0h/r
9FkGOPaP/JBh0W+nVlRGOHO7KVlshfjO4Qs21rBQ6LRppjlU9A2yOH3iBclK5uGXDWLtu1FbfU+F
H/NiMTbs6B1Td3HvkPqxrJOlyIWTyZ8fIhfKSRmoCWjEIj8Kl1DGWnQRkPIvEwbYSFlxGAkXmxMd
ywh0BWFIHZUEUKwkyOx74rkOiK93tU2YDbO9cxwdrOUQBr6zdJ8GtIge8qLh2MKsNaNitzApFDpd
U6kOY0l5OLxlzZbRD/ziSMoQ8ltJcv3bnneOMtwuLZ5vlNTaXHo0lDwoHQ4wOaQEgRLvYvk+xyHd
q2v0Wk1ia1SrfIQvWiyyN01Yw9nD4jaKj/XUMbxFCb2FTTwwqWbHDR7886yQNFjrmaBhhW11Kwzd
TbwKbvQPL/zFKskENH/PlBjnhaR1E+irYYwxjt7rESlMP6H2wmIFkTHDCMvow03QxpPaM5CYqkVN
Fz4kHymzTAhbq8ZBd6bmDrZnV158Rr6RjAV+p17tlxQlZTNWHwB9s1dpUQxl45R8xDziY74rF4/J
eJ+KfEEoVsZQCMoJTjwyi3WxyDC54S/thkOmYyxcby0wFZn6vG+fpF6SIstxmWuYM3c6rTdAsOaa
J7fVsELU7oTgKgZ0YgTROwkYtUF2dnqfJn6b5yfikGHxLCUYaHP9Y9VyXilcuvuw+mJsZ4AX6KtB
PpYMQ7JajCBkJYo/1G8Uss8+Po2nPcAfs+NLLS2nR65kkgU5la2vfosgQFlwtcuWJSbdAmjKGHII
OUeftzwur5ks/C7Ga4Ayxj4te8t/UnIaXPfFZGKbyWkG9GB3Fcj4l5i68YpJTKr3XwO3JG54Nhol
FLYmQorcbxZsCUqsI61FhKI/9j5XjaEqtOE/woftHTImGE+9G5oBIYHqQjO1enD5gyO/0oZoE4nM
3b79ySAtTRe5QD9/fOyXNjMl0tAwJLhf5CrUzij9wrYWJFlOqCY+WYIypsxQWNoEEp5ypNp7Mlg3
6nO9P1G2B5gvZVti7CBtkzDePxSpTkXuFw5XY07Z1Oyi4X5qiiBSfK1AbixXodIEtTqVhDV1QLqk
C/KlJb8Rs4eFqUin4f+m/MpeQdd3MPtLpyctgvcn+2AJCTcX9Mi8KUYzMZGCHQhw5m02Yvi3o/8Y
Kt7gwZgFkp1WT1CAXGQWaJKzKS7bI1BT2/GLEhQsFcRqFDDf9lUCftlD2snZZVdaqfeoack638YE
NX3nXac3w4dszWIQx3Sm4NzcozBm1DYTXexFleLAdV+uulLMUQXxpC12wi/eqJD+fspQcgXE7gqz
gOqlFzkhyK6eR7kbYDBr6b03psHdHga7bQJK+D6IKMtMJLYuNy6LeWD75NvZPTxvgVr18y3h5IpX
qy4T90okzVDIF9/d5RJ6/ado3QPrbELYHBBfvmod/XESOA/uh1TGJouguAX6fCm7VHuenXsCSlxM
L/3bsVmG+2lzSL2mkvTQFG94yJpvdmswORR1N9hhZvYxYmwm5ZXTZb/0ULkjCtCqobs6LmC1KW51
VAj7qAB8kdqjfkRpp+sMDtM9+XTZZypSq8EWRNCCFuNm9kMJdap/zSIWLXIYvox5RcB0FT15llPk
CTrDXoGRpQQ2xGmIOUYFIefM35Jya2/qmbQYq0z27c1PnvOBonyq1hnsU6pQuO1VlLK1O4+2Plq+
yK18HWzVnDKN2lMIx9xUqMSwCeNd3nAC8jvJivRYHHDqdlAQDo7kBmNdDtxr/49G0bSQ7PoGNWgQ
zEO5NrYOcx19Q8oFt/znJSxUeoqA7ORRqzE8JdRH0oGleQMY0ffqyrxEgLXzquszAoA/6JVB8XLV
Q5GuGkk9z1r6WhPjKQybV6nB/go/L38VoTlHrja9u9mhCbxOJwinvaoKWzqEsdskpOVgvtBsk1yc
U93kmfa7Wi/yvOf9a4v2uNP+9UbOeDPTqdahmtvsL2vk5kWhFrUsQc54b36DR1uj/mjyI2aqNeM3
bou0UXF5jR/lGtTqONE07ZGMve7vsulcnGVYASlWnfcvDFp4lWB+18+AsgEY8Kz1es7qXvTIQSHF
lvUMv6Vsgycuans/CKQFgx0+q2LMdVKKmslskap2nFsAMzD8j1T3Bq17CPmMYEes51AYxRmdXn0y
O1uNEg5xLEV6y00fLv/Q1ClAf1vRTKtlwUBDYEPWLxyk4SjFn24hPkBRBUPkQecBquBVhfmow0KE
sfdkVrOJHpjm+w29qyQnkdgBWQAblPBOwv+hMaKabQmFjAr69aJhpU9pLZXUE5F7bWjR4GUZVK1j
cXY8Gy0um5s2xK5mQ1eBqSEbKOI2uZ05qnZILglteplCUi4uVrEzIqeHEQYcH0/0WfQWdJaYSrRZ
NQtkGxc3td4RHQx7IR7ONA4xwK3c8CsAdJt13EmFhS9wK7RO8B4mqH4qOrUvDa0mmzCdLgRMdNHq
DlsjANMrujjW+F7ckcI428EoyaG4TfcIQR3kOaujR7+hsJblVBmgsG/jO+3GaOvw5WGlz3bHu6Wm
ZuBSdtQ04NK2TEBWXrlPB3MHEIlEIS3nxVTBPEzZkNRgYKhimJ2BE8T1eDFkcu8Z5EX9HVuk7l8T
7b/Pgp1I0BCebG0A97GoJlmScNlFwAxw8eOhNUqaweapIWuzFPaoilybNxLZhUaFEthS3E/ASley
Bx0ivwW3dY8cGXKUS/q/uUsxegHZhewGZ8n3A9bwgycbnDDaTAKn6Qh/BmSzP6Ssg5373kqQ/ysW
7w4Ae5zlqgenxC2h2CKbCXys2dR5oHhskLFUNd/tIAzbunxpozQry3DvQaSKkafATT+KtnTh8g6Z
MH7lACBTqTt8f5A8jGaOoNx/uFHL91qhN6lzCuOLmsgaWAIS+c2X3tTN8ZyPXD9SXYWVv9aQX1vq
YZ8ADLeu7kiaLtLu/uThp7U48j+hk67OFPIWziZAu2UXxIpub2CJKqALcGlfTYAR2IFDbOD3QBpP
c1OAmUmpAlunaPPN0Ch+vIQ/nJLROznX40TMNEeQaFmhqeOVaXmk5a7aKrWPwrdwrORbfzIRI120
HQok3VM4T+U8frHugL4WKHd0v+1hWaEgZI+10dc3pqKXSdxjWBuG5KsS1m3QTU6EEsvK1M0E00gY
LkaxqBsKuFnkjKcm8NKkRhmX1URRKZWlhJAh7jv2zB9Zd7ukPKhnndCw/E9q5dl4GlIb2AQzdyaI
eqFhc7Ry52JQ4SWDFp5IZITGNbip585XxUkrsL4pfJARm4SaZ5cA67SNJ/G4x4Kv8JWdV9ZXcqOp
63Xjv+mSffPziV8rAgncs6cvAPN2165YdR0Z9EmYxrHBASU8+eZvEHibIblJhX9/DaLOo3nzqabq
tqrutQUirayNZzwEMHrA9TwIipfA/6cTw7ab7SzjLL6/XfElV92oYuRAibOcPnbXQUMVh+p8RIUD
zcDGbZtCHn+Lc/DE2EkfZSEIaLh7F47Y7T6Pq4Hh0JFYVXgpqxYcmKdVipu/PJc32yuWjYp+wUiC
7dy+ahJ1brtkedc8hfzL/RG+qjr11264RFx3syG+JACYEykaN116dxLd2q1sk+q5G27ZzCXkYzuS
f3wyHfk1lxKrNqtpNsP/At/jL+hwnhtVDdc6LM4PbrF5EYuAF/WD48qr72aomaIhxsN4412+lV/g
AWQuAIpzCls1rZ+81x++WeitMtXXRrRm9bTRvDNv86kz8BMoexZ1spxswNIIsTTnuP3eZxsKxDsr
qfI3MoC6rwndtxOkPBjmt/BtGK1pc3SB4wYislat64qw84OgNNQcPPoKTkLee/HFpsqWJb1tUTbg
zZ4jNYBDkJ4+i93Ivp8Kcy617hilvPXa5rMRo8gE0cvBXrSKvgY9KqZvBb7XfDoV8nNDoR+u29gq
gtTx+NpApQ2y7JRGe+oLWtDM6PJF1K11eqtREH0qOHLPuzjGBCp3O5GafTAlupTrO9jiA4WnzKMC
qW5uoZY2xwzfGpOkwKmN7BoYIJDpfBm7614xb0A6xpJAMRTSuNWDJBnxZoayd2414Aps+jqNY0ME
LB1416vZ0j6K+mykmZNs/O9AAcq5BU60kG6aEtJ5sYIS3WAQCDW51tiWWzPY9gAxHCBVDU6NupPS
vHwxcMxWafonO2P9ixSXzZjIWA4OvjdiboPm6s7p4YsrzKSSHNutoHfINCKfOu/MhK+z7q7wye8A
pb8nsSzSacrwDW5j/2RixtCPpZE5oT46p7Gdyw8uVcvniZe6s75trNniYJkt9MvFt4YHhjVJ9iPS
6sxMJBcKI27onccqQ/qH+HcyajBk3Zojg0bFB88YHJYXpbbl9Ivb0eGNrKWwodMsb6G+rpeFdTNE
VOyFP1Th+a2ry+BCWdYk74zpuHeHgOi1VjOMhb47eVAzr55dHCCSwyMpC53/+mkLKWP/sSaMo6Cy
rI18jMMZW6G5hzRX4XbIvFln2uodVzlxCAz3mcU2a/7ijYkLvPafMAFpV+MnCgxoilQXoOUFM+I1
F7iiZlfxtqPSFZjMj7/k5ki0mJUgJRFNwnpkzAmqtFSrcymjjUmmz7uu5Zwur0B9mN/fjUMbidhz
9kxuTYHGWYEyzj7WNzMOXxj8WGkGGNG+4tvBcmKk+pTH3g3Ah/yjnEKTYItF9OXyuFv56eGzFNKc
jnf02TNBw6vSO7KibnFlrgt+AZwq6TyfD2iKJIOXMqYC8KoznLffClX4r09MyC+qmnWsMTihWUCo
qhOFPsJL6ff4tb4QrptMmdRPt4LBKRWSfAvP65YGGpOUrSNeZtEEeLZ9fzeyXauBqSfcBU+7j+dH
WlJ6YRb/2HiqGHW/8UYZAStyJPaW/a1r63RZNXflet+JAiK9JMMSv2kLshy+qGvqSPUU6+Ap417h
8CFE0o6TasBIV2+QsNfIbWUypGGYxfYo7usP2ts4KkDRcZb+xEj3X2j7oqjdtJd6B12P6YEhyk4w
VbEYMD4Z4BdI8kEE6fVYxBlLkWbAJAnOBRwocH4EnGD2dEYHWdMiYZb5yt1SOIpQ1tcIlPFR/D7R
978KzzMADNYUboqRMJLlIHygkjQnyrLEkkx5J70TxQZzjKirWiuyPwiHNOtG5D9u5J35LKXa7oth
3go49VuM5FgMB1t0sfS23HEZQO2I/dC166c3UppzD3054OIIHQCXBmtYGRQBuj+zsQgB7CYcaeIg
JGOaXfZBZJ7ASicjxBKT1me0bROMt6558e7wU21bfOc8b0y4w8IZXldrD/xmABsZ1jqHGvj77rbH
DbT6qv8CryD8qdk7ygjql0yuDnqDvEtMhS5/kplVEkXLMFoN2k0s7tdiKX1YP9phc2ZjqndIYIlz
1WFhD1eKoCKwE9hwPPQFZyUqryxoG0fKyA4/4QAeG3Zn9IE7vTqby4rMni18nq0kouEHmHA4+FkH
3oDyeU4u8xL1o1u2e+RMXpHSK8NHgcZMFqZk893ZOl2sgJqa8lR944h/fHJ/9LXwddAwgcADOX49
yFht51P8QbuHZpZe7ZJr1GFMQoG9aSh/IwyI7uuSwSCst/3qwW1nzyMMznewFaTV+42TwSr/+qRg
5OwSLjqYo4cbVhVmTOjrTkKWodDkXWc7V4U+Bb0BjjGecpU2Fhyn3lwo5wSl8Jjhkn8h2WhgJkkJ
QvXXBW/keheiFWPMsjFDxyOEydQTEypFLRje0heIOwnqTYlvdqma3Mug0J7yUpjH5cDqqwYwNO1r
e75YL2IYhb2UC1d0PdUVTW0Au5hOuzhrQLmZDTE+Ij7kG4lnuxd/GcQKhe+Oi3jElNp+4yuzTpBB
vCVcoZUhIeYRdu0aSOtpuFGB5a2QVuICM+uMHEIy+dORPSQmI4IyZAj3uuL7qD2ATP0yiSiIS4+w
isQkicrbB+0mdnvILt5gS1Nk7lalpEzYxWLncHKsvZqKciUQYS3H2JLNjNgT8+cYJOtC1e88BEHg
ypTfLA0iIlUw1qvRi7WEhR/vKcSI9zbMyYZSc8YT+zmBFsuXYSyxte5D8XqrHwfcdwIL7Oaiz2aZ
JuXxPmMpi0WiKiSETSTJRga57scgNrpIxMu5alkaKybYL9oI9EUC8OrIWMBYpy3iVEYp8B6Bk9cp
G/8y/MqKSmD6tgiK+E+aMH+MePZS8SqZHKS1Vbi9yaaiJnVnwXodmpa0dhz92zQgu+QB+TaJfLSy
uCMXFC7oJauIcmL+2tChR7uLFhIuRNou61lNOxgB63/YsLWsjHrdwd3oe3OZAHRHeJnsyZdGW6pv
ek12JAedZuoPS1tm5/Pwhy4+l93GZGXRA+EwQbMjaKpepGzxKhlRWnFKr7X3uIFaTBY59RzlY2gL
s308J5ghWd6/2PN86YMK2uPY3vReZuEPLmTaeSxK5yOgkPmgxh7Ln3XmRKgwi4VYrIL5fa4kWP+k
/1pyj7HnooTl3vdCDe83Av6qDKx3NgpgMg9w+J3OHm2yX6HQA4B1PbOcExdThWwk0pMbxp8Bkoec
MObrqW7XO4fgwdzsTzkDU1QMUUhKdhL4iMAIrq2tQ3NAynfklh2bXDVCLtTxNLjjNn5FTyNHUFUZ
aoIzCVgJY+wY8/C685qrv1z5xt4cIyeIgkTEkTGiF1wWf32E9TKMjJj+KW/BQC/mThr42sl0JKOn
dqtDxN70LqucVMVkBwfYyAIL61WRqRfXgobozvhesXHc+f4XZeFSzDVz7cvctJzveaWq3tNaSFJO
lV13hTO8bfacBzxlpM6NcMkNsaj5/8ml90WvE9gw0IaZemN0vb6ct9M+B+BgS4Okk5Yv1oMTsrX4
SajnbjJ61068tcs95JGBuZrpkjRB8fdNjKN2jmsGYV/3ao+ZmmtY/nY5pKsgF+JHygQm6uhzlmd0
ApOoTlbIx9hnxHlLvzRVxcKfOyFNr7PZpprf2A6D4l7iLwZipELOpmz/OfRmpTrlE3ynY8EHZ6VJ
Tq7eMV0lBfDDt3c2gpXWfFxqLfqX39KZr+LVXkSBuvk+hmy8EGza5zl51jn+QUSNgJ0GLDnLWZLO
giIQi2dSpPYsML7gq6L2xRiSMfgXPnraQRk4IUXXEQxT8MQNjPIvpPJpE7owWBg4nVwz93d9TF3Z
AtOUk+p92Lmk6r20P2DEGE5qFUaWVqyqlfq7OvbEtWFAxgEfd/wUvFhWNK2ZCRuhJIGpLHVgjtIq
3YdF8NDaN36rUb7C2METa4gampGT1+nfnN3xe/be+UKHdYTmoKUZqMtHcl4hQOQuREDXNBj2imhP
9LGhLjwgExE6nuG5IACW4ukPytXq3VXSAR2eJKszCf9MDawCoSDRJ/6HZ3SmLg2k1j2If3EORxEW
CKqYl5J4ZiMRSBSWtelM3e7JWwCgiDc2OofX5QF7emoilzPJQ/g6o1Mg157Z7bPcyqcqEGiRYECT
iaSQ0pB1bCgn7Uk8FGQhEuoUkh6jtrH2ZOey2kE4xMCQMyxu7m83SaECEMoQbmcEH3tO5AFhpEI+
H1RqE4XHTLstF0z0HdfId3mxK98eR0CwosTqhVW8NkbFt7ZcRJbDfIzrx73wWJscYNhguWttE8kM
Pmq6r33A2QtEF5FIt/bHxOFNhb6YtmIbZLhA9AwaPu6rojOp4Dv4fC4fynwI2d7h4NxI7Brg0w/y
/6sDCOAbIAXd9tKc3Wc54Z2Qwwf0p5aiVx1cKgmKk/x28wCCLi18O+D7WpSamj4maksHsnpaP9Q4
W8TFJjk+JvoRsp9js9TcZUvGy9G4Gpj+h/jN7MgeN4jZrwaVvBg/OZf5RPvXsALp6S+k6N307QqD
e5lGH/IuvKTWCooj/BvLLjwcThCrohoHPdc7lML+LsNZ4DQjVhNa+T3V7+9eNPggXxH5jjQyYa4Q
m4eMNRDmxbTIJrgaTNAacsNWAfY2lwLX/ccH0vyZft5oMVtxnLWyEFkAzUDscRbekro3P/faBr/E
ctv16dp3SSrhqVjf4cSQ14JhvJVUnq1S6kBLDBKVqaoxIVmDqlN2vv778ArZkoVzfhedUeK/lhOU
ShAZS28naK8SBUhKLb5ixIIUiosAyc/8U+p2QSlvSwyQWtbuVkTUrPU4+5Cme5fH0PlDDVkwS82T
2hLcc0HWz/HvunwDEyHeALacsGGX6VR9fGmGGAbiOyyduN2P7pgiJ7dm8ONu0N4KNmj7OCAwLQrL
1XmLD6eFqgOHF2uqUVuXisgyJzzdxn7phFj6tKNNwrtBJKJFl1bFqodwcy0Kv0b4yPbAt0qKGluB
yrYT5vyCAxHlna5Aoy3xUmRGOeOjRzHAkqi2Jc9JAlOc1mknIxfg9FdfjpReU7vFfhzoew01fQGx
nHOFn+dZVht0rGdYUlau8A/EFArCP68J/+f5zmykQjE8qCTMY5YcqRvPZI+Z4iRCxrQeBdQxkNME
nhuyrHEao5JL1i610jGWW8TJz2eduquGqY/8szfNXPkabH/NogOPXV6TvR6YLLiWFfFM3EZHWzXG
TPHhJ+MLy47JivCOCEmZwgdhjN67O0hclffQ03PKNK2ZnJHMljFYKpTk9gd4jVFD7fWvta5DJRWQ
bl0DChaaIRgtbLwzDXzi+21wbfFKxbBKGepvUc4roe36VdK/a1UbxST5GOXza7Llbp4aUhlx8DC1
YGCh1s4NnDPAa3MJ8tW6ejr1xgdbwgvrk9ArjLVxgcLcj3aDLwcvnWF+ecmuFkVuo2XfyaoaFzH+
TwNbxz057a65ALKaRaRKfxt9GIdQ6idccO7bMlqHY2j226Q4wniFhjeIuBzsqhnqIluLkTTj/o5I
AMRJWZO55Y20OwUnsm6HYWJHi3OS3HeZvBIERRFaqTjJYJGkzWcLW6iPnwbRAlbQXRxJeEzlmgiq
RlOtVGOwYee8A+hKule2qECXRnjM8v/opL2tn0YYhjGDbn9rKYXhMMbZ32X6pBfnuxhaLIqs4h1c
mSjLzKoVpsC6r0ZXbx9TnKtTG92fDTw1YKb1UBclZt/NIA6eRdCrVWBxA5pIiXZ5Q4Dg4udgru7H
uDr9wGWwzSpLeMsDohU0/FvDhdEXT//rjrLdZHXDjcx/JRTW88Fpf7vZ74B/6GZ0dHkzFq+3QPQH
2DXtQpLK2hYaRzjNlWAzZdiOBTGt15UMFfLrOzrrO8evnnQi6C+DSogT5EBbKS4WLwdhbPfzhZ7X
ciNOgVSeVINe1Eidvhs1c4/fHLnQxN1x8P9X5Me4PYiGvfXc/MAHq0Z+jDJV8npR7vABeW9bUL9J
sbK1f0ihnWDpj/xFQiER3Y0UomwzDw/F7Zi0ROc4gBUFHOIcDdmYYTzHz2JCbEmUt4fdiCeBploI
slbRkzAp9TBXgvMdzCHa7EWBOWN0mni3jko0QZQZQGxU9h9nhIR6NO1RfxtQip3IOXdz1BzRe4ai
d6+0jkhjzo6dJ8I6pwu2Hhk/QS12sv6C2obt/Qv8mrdx1nRlyaGnvXmdk3IZSgq9wQBRbH9fC+Bz
GDOmGCZ12UhhM7lBV/z/lluAe6svjpuKu/5126HqR62gj3V+dZ3L3SXSBSPUCdLEjQsqd6/IbLGS
0Bwf+3qBuMvra4srhcP61iXt3bLZldHmjtL5Cn9BFb+vjKFZ8qslVBg4T9kKkeAIfKNNcUfuixGP
SB1+YZ7auRojPoOEOm5WqZnaANPC+l+iPYH0iuPUH+E9fXC36qNue8xwYG2k6uccTA35GVT6AmhL
ha1qab6JiiOzUiSUSDG9PfWDXpUL5fXod6xSXRqh8F17gtgjfixqVTdM9YuqzqWBbqkjlMZHTJso
5eRAkThKLk5FESf/MTL8CgjLyvZj8iBwz2AOVydqWXJVigDDA/zaiLmv+pBjwKtijZvPmQP/A/Qa
Q9L3tcZORc25Emr5IGlh/H5HlrJYFaPgN9XZMGilXhBxrJOL8NVtgcyguFSawUcWtaxbUGMid857
TCbOQalcxJu9XfVBWCMEcmWXVLQgaCVKqs2ihao2skM2B3z67Q3V/Ydpun2Q1vn+meOpnP2/3RTN
JxhSsDZMO2P1TJ+yxtHAh+yBIMkrEOtC3xm+YTneIkkkuaW2CWPto0lL1UbDLm7nxEQlF1m3k5Wu
9w3dIB157Ny9WO5MmIpfOhKkqdavCk7njg9yENgAhN3mfpUfIYMYsTwiXD7WXGbY280z0jfItC4g
p8ls2dbgkB76PdUFzR2EzcpTqzWJxHAwEEk4FVhn+Wy7S7vQZjpOcXrjz7hk29CTzci+U5ghFWV+
zL8Qdl0w0gxJi/xfqtyy+IYhOOuJV5w57Ysspgf5V0ZxZDUB47CwXX83ojom2slRB+g3XDKplRQS
3+JzPSao7yotKjJGhs6GOupEW0NXCG2DAQCaVVqs52dixkV01C4HFPI2Ibj9iuy9yFDMbcYx/Cr5
xhJa4OM92Mly380rjPbvw1pwbxpIDOE9cGtwlu8xo7Z/WvCNVM4tPo6crRtYUSC+JmPygmFL/sJG
8XYRxSaaYIC1v5xnDowviax6zOYnnQVxCOsLQXEpCbpqohVphTux+h4WoGpqaQ7B3bqZlwopnYYX
lsKBSoN4NMKdS/rOjidVdM2/1exx41talcsBjd1qR3NDC5CHzfzI6Q8oNWr0jGD3pS5Ad5ljyXC9
24uzBgM4CP85mogqZS6t3KltXBKdX+N3vnKCTci/lm+tKmcpLNped6JRAWPABi2OcJFVhajZYK29
melQHfMrSgNv7KHOYU3Ik+/bhs8n+AR56Vq3grV2cHXCUIcm37sKIc5Ho1qDcKD8kguRjt5tx1cj
oIAwRCKXAon9A/VekLSC65dghGVdfc0KNTy+gT+LaC46MycSsKZD6BN3w7lC+AfOphWxxEvrREvs
60VE8vqJq6ANRcKsSxKN5jIZlulAYa3EK7W/cGqqSZHRIJQRwq/zL1aAPykW3NPy6DOmikTjDtWT
QwmdE9Fewb6W8zsBJbq2nxeCd9xNQOVKSVVkmpT2iebBKEBoMxn6BmJKQt1dPR/uD/IgZDoZoN13
q6cq1mctYtabbZjeIE2GhuhjuGvIRyvO/arsM2CWru10ODTfpzGL2nfz3UXpwKnbVgpxLJigr7tm
9UJs26ZMlamPSIaPpW+e1ntADw8LVFvPrJJB3kwFHfLZyBUL6Jh2dzriq2E1vdfklZEMX8elwzmd
5a8oRauRq9PqAgTPtdIdoreh2n+vDfE97TIvm3bM1I48H9FZlsvlPBs6d+BsXqce8GQmy6P4kY7Q
4Zd8RkJXflalRFa6xrplKxeWM+WI4Rry1SG7Mlka1v2w8zcX5z7bSe+FA27JpklyaRocU39F8FvB
5qGeK6jiQKlCbGYUKFARem578PBG+IyjrcVmlDvo+QhKKfDV6AKhjQ0nl0JjnQEbHigxPUfGYbGC
KGCiO8Q/BT/8sTsNRk5fQkFFVZfutQkXZRAxdUFU1ETYo4VG50yYIbG4IMVNiuF4aNYNqS+4cR/g
v2MZDKp/rL161wvhn6zTi9BH6+ldrsZy5nkBglnfv6I1K150swgnEIGWeOPsnnIGHHRWuYi5ck+q
Zb8HxJumNL3pNai2dKeZ3u1AINCbf07bff4wBwK91+YApoiH1HLx/n/CjlIlWdvp3VWTSKRJgRBJ
rmY12x59B2NiyNr7e3VyNSEGA9NNGMfmL7Lo0p7zxqYNciKphjlC1jOaa782Vq3Vvb48zFzj5icH
W+rBwZEkAyn6iEzI9gLZjy6mw1Q0mE9aReB43w6erf//yHlGBvMebwGkqcKJrWMiM584zd1nSrLe
UyIAO72sRCaF+s+H2/EQgXfR5YL/x746C7fOY1N4uSdkUT9aZhm+65F+VK2qh3YtF4A4jdo0IKc8
F87uQ/QeEH9EfuwtHaBfVWCZhwjjbeSLQgqeKC/mn09nb3EGdZBuYQzth5v/3NxTXAjjU1pa7LfI
hfvOMhohdJCk1PfpbDMasJ2N2OTDdmECq0xV8rjfgxy3aVdLLpWhe5dWp7Rr+npiImT215AJf+x1
4oouzWIZ4MmNoP/DQ4wI5d1SI+LKL1k0MX3nQzinOJPkegBStsKbAaHxHiSzQnn4LYX8ATlsjKeC
SXWWNqJBjirJl59gqkf+WuaTxqovg7HSanBmpHZgQCol1v7vAOlBI3HnVMAYKnYnA8NRmG5pQmKV
4UV0DBu8jIVtVrgMUUTmbdVbpahKuRRdKrWjzJVxmfESo53hNj1YYR5v6XJucuWphiPekHaW/tmf
YmwSxeZTfQN4CorMzNMSaPxcNYQd2WkeaY6RTGQiSGIOMC5Wm3FpfuMStR0uS9Eycqb4MLhdrRBs
H1rulsIoOnBnhoc+/5sKsZ8Isu1TzXyWX/jO942nEoTH8EFPg67uTROeb5QWgeTBIaWtxD7EzqKK
SLmYZ75qV22vSXBldjYFgxUm95Xmg4WvIFaAwFqiERfnaBvr2JUWWAJxiwAlu/MpYkxDd/68YFsF
sGpU69VDoBREVU5gwWEkyRdukvUrIz8dBHGQ76mFLbSVDICFp8G1lQqYbZLRJ1b1SJrOQ33Y6plB
6+KqVO5wGfdWESQyIew6PWaWpuvLDuiRHUjH+9l1fSUyfuJBeqIZSgnlcfnFWPQfOxGWBnGRx/TA
2uwnEa266nn8nb9kmr7Dfgb223MtklQq2vfoVlL7VcMAo1qZ9nkG7qkQd4oKNmv6LF/ym4+xeTae
MsA/bbTf0dqUWWhd6+tkrtagTKXfhyJkj0vIxieFQh84By4mjwEEH6M+x8Y6DkZJEzUUIEa8K/GI
uGvcLU12ppwZJ+q34FAQxe4dJBMTCnSuIWz2nDhLmU18I4TQanbZ9i0STG7gNxV8GrRkJ1OrBSAY
/ku0BAAvVkvSLu9d7fr36Kv5FRRJrP/PiKm4LAdeJjEZ1hrUZP8eQj/AKsW9zIc5YU9qHmM22iUz
ohiymaMeaIl9Rx/e6I+0E+9HBtoSI05x1XYkZQRpL+GFaitAgw10vsi2oBfFj8WWfuipv94r+6Tq
FFO2/PJzwIFC9I9Uaz3BWv9ElppcCWxXnZb9XkPbfEINlwCsaVmI7jXcyLPY/ZSx7Oe1XKiKR8kk
7ZpljHrqMuJxoMs2PhbVVIhV6qpCzGWxxF5DSBDK+7x6u81ep4uzrmkZN3Kti1kryCToTOUuJ/WH
bjSVonID4h6MkXx47JGJXr5C23qv3luDlMRiFsUKsZikQq0qy9WfD25Bgz2RjE2EVPSBZ1HpGcQd
ZNSbql3TEnPJvfTZlhNGd0zqzwHJeK9wgIs0gDWFhJ6aJr7Uwf2OSD9V4SJZxYLoaUEwY/BgKqCt
qSXBvs/fetiI2XN0iEpj4WpWkxMLlwdwzZQnFms/gHWHTTtkmgZ2/g0IaNRhBMQzgzRQL9o9jbZo
cD3sBUBmmM7cYAt8KrDdL03EVXPNjmlWSky1cA1YvZ8dNDB6ZC/Legoat63/trfy2TGQFDD6zguc
XbipYzBnbVKQAHwj3F2WtMJPCvHKfrE/3ldxlFsAVBqWuw2lPsxXdbaygWYNuBPjPoCgvnnUYVZZ
EF/r6ZjDt7pWduSu2xwDNS/3116Dsdc5jrcNxiP9YWBKge8JUTPA4lB0X63N3/qGE+A3AlF5o6FG
Mz2eUrrSQcuTQry1xMf5Fi2QFn31T/pfQA0lrvLQfZyjP72ECu7H5yTjdINNPdFn7dtR17wo4FqE
YIro9SkSNTI/EdFSulpUmajZHnf2Sv2RDGL1LCByag4SVJlLdrJFMtY+VZR0hOPqIs6niip1z8/R
opKZInH/pyN0uJ8ovUd7tBTvQc6ul6eXbHf5aI+xT/HNjxzf0iZziVJTER+IBIUuCS64vwSSQ/0w
ayDQk1+BqY0he68rRUwW759MW11L8Kvq25gfoKxVv+wwPeMheH4/pord7wcY02JlFqkTn7qvP3BD
Ksj/PDThspf17HOXOgE15q7xc4MVKft8MG0CwVeg8uGgK0NBqaOx6LwmPpv1a6IkPO1fV0ZFW2wZ
WDIT4SRyAZ61LMKrTFZcO/PLRmqbTpR/HGQZFqIGnlBwl1PJtFXUhw0+0NzpUzaCDQUKZbOWtp3x
6lS0TsezuP5h55zc5aCVAEGWkUgTdHmRVk/1t0qtt4iBOE8zA1w9kr6qOQS9vOled6ILxhSftLO+
ojEEt48qlqahvgQVqTaTKnzPOyTymlLfDdFvII0rbiQSQfXapbRFwU4taxp5NjrbcJ8MuSfAOTb4
jWYO8YCD028Tk2UE4htkrV8wZuLXdZ9kQGQZIz9eSnNmroCX+4hZWYa3RGW3b2ac5Cdnje2sFliT
UT7Lb4se+XCTyM5ZWIqFjVBfA/j0pZGFcgUrcSw7PzoXkVqiLMo7a7bKLjE8nc+58D93ecxlAnaY
sWlu/klo0qAVdRpblHmlQgcC7yYgMU5UjaQ9KJnyddNWPQggJxQldcxM79NDSrupiL5cHESxHjQh
zsktlgr6se5dMnpt3SJSPIvP0KlsOvMe7T+lJzxh6LHOMtGn5/voC1XNFzVd0xY9e0UZRodBwNZX
bK7ztRe4/Iywudeb2sob5f9YoW+bCw2p0DP0AtQDYtv6iA/ixyrFBJE6dZRv9aaiSW5HTqA2vvdg
IHmKVOFpANScYqKSoaxfy/CUXunkWJbpD32RYPHfryOGOhwOEPDk8IOhJXrirOu4ROJ4oxTjHDal
xWaB+21s/e9J/cbN3vMVE8dbxqSNzSQ2KbirPU+QY7kJOo8dlqI8XyPpbWrlm3VIlFasE9dUFXFv
BB8nDVhS3gpsf9NDRjB3a9trvRQd2MwCclXk2nBCJfYUR3QyCkieci+DGtFlT+H0gWuP8Sp+013O
gVeEczr/ITHKBmmJiwPRd6TOL4W32bjBqyKBEw6M1txzmtzC0Q7B6OXRn9wRAKxw/Qi9zvrZu7t2
Wag9psIcRPyPeOOSkKsmFLz09SDlwuoV3BIcz/UPB8R+Lx4esRxY5qyAIFwv0G3xAW6/kUorV/e9
ab9gZawgXF5iM5vZaJlfCmfjun3bl5OARVKNsKMTzbg5aEXKTkRoJwln7EwhcRMOJCfZycxJ5HWZ
0SEYR5MNwVvV0tQS/os4Rb8bAdhAL24A9HQUyh9exxF/T4mEf0ks1/AjHrDu2o7V3qyMvtLZHCfx
mVsZoCmxAxfnnnTupwnaC9NdpK1j1ctLemUPDqTavxwJahJnt4R0epuOnrX27M7qnWTnUego27Vr
7DJKfNjthMTxnlhUCeRiD8oJ53o1rbZoHAytx4iVbtvBdomA+PmgYf2OCBP5vUNF/t3EMXLSkxJg
QzIloJPU1A5oGrmNphWw3+tOyxMWf9Fp1/+aPSG0LTFVYckzjlTLnu+pWW0rYHagr2tXiixqY8SC
g1c5Y7S+hwLVQu9wGQ3tsbdhhQ53IKJYtnxteQ1FqmRfu7GEvm66cZj8I5ZSHpEgAzA0vOB5j1iA
s/p84H8RqhcJS8CDyMFwfAt4mCnkOZPVrIA5+HtXxZ+yOvolTdbJ5L6nSfaWOTpjyxDokPI6oBGF
KmHGFs9ZK+EnOyRWI7dULx3mjSjswl2bcnyFAqsRiNzYiBpkxP+RR3DrA0lBskXgpLavfFASgH5P
Jorl31BKvInycvOGraxcm4G9zrOWyF3acD0/ecZppqSPQOIV+wjbNBTccM45qN7aUwsfZq36WslR
/+x+c/bE0JLPW7TtVDQXNd1m2Da1mGxcxT1icv/rUz1s0N2VAjpGaUlfGY+qKDvwIRsSXnpQb1r0
k/ieQkgvvh/xCtC2xO1MGoDOyhq+M+UzqNDE180kAKTDdLVBK9/qkmd5jQPxEBp88G8oG8wVr42n
WZzwlZsltRJwIqI14MqYrlwJfXwwzWmf3Psrd6yaEDODDXNe97+2gHWryCqpDA6z96GKiuuUCGji
cdl8eJ8iy3Yp88uYarMdd4LLMDTYI8KQPcusFh9ktKcW7OTstCxGbzcbuNlSwZcYsPnGoZ0fchoL
RvpGSoXy4atp+6/gkCJDWvndm6+utBn97PjJEmP8vOmsnbkLDaG2kRoa6phBcoXNdSpmkqKrALh5
pGlvqkdFFvveputHq3LqcZCO1zNsU5wQUYsYNvyYpDFMVWFJp7ZqW+JdjjQ0ANzTj4pdSpjoaibD
P5KvukALTN1Ks2Ih8n2HUtp3Cws58dxvdqHDOac1O6nVSvMl5pfiO2W/myX5yxoQZpSRyeHxkOVs
yL7yhP5s6EnCkdZn5awTmWtjp12sJkA1+eUklVnkdsRj/ozy1zVdXiA9s1E+xJEvN2eBujo6otiM
46PyzhHd3jyavm66DsyHEPTZgBvUq9ftyi3iATulNPw5+mwLJpamKZE8kj54TUsbfBXKXkUxVBd5
RJOUlTXW1RV4OvlalsbpvSqOW4uDEQZc2B7Z88ZImjRTc6zNLGAz6L9MaMCwjQftaubvCxNfnuMu
z2UJJbj8x20XfVBU/xjYJ2FoETVWpzYiaT1okTCNhcjLk1xKdohCw3cetR/avaTK8MXRyF7Jzd5L
YECC+SJCJDf0fz+Q+rM+2Mkzmz0UTyCjUbXUDrObgXv+WKH7wbvo0SVBA9VdcjRgxRhlE9KqYXnV
JcNDUDscvNEXWaPSyHBg249mF+rJcPf+/JsEA05BzzkLViRHoqZu22Isdm6vJnyOeXwuFJ5huDuJ
Dbmc8L8GkxZCRO9CgbDdMTdQ0QhYu6mCQm9NAGbbIOTaObWxo7K/qzQxckvME6laC5vfHSX2ebw8
CAjePCs7mbGpGLtkcAeJBSkN2Ho2hL7mIUckAvL6zdVbUIXFP6HnxusG2GDQ9GhEYFm953CDhQ2W
1sws7ncyo4HCh1CRBNA0qr6Sjx2WCzspdPynsvwE8qWU5dDy4RiOj+iFR1vfhlP0kzo5X1cI033H
Rizo65+Rb/cvV5+4Pv/RVjL0eQg7/jCoO9fhVinWL5FrIHIX7mk6h95qjLl6Ur5wOy+Lgi0FWIAT
8fM4GxQXpzRsspVy6GdysHfy0ZNRS5+VBQYSLoWhe5LlGsRyraJ32pUH6365eHZKEn1wfNvIOyX9
Sr4NUB0mfbABMuMoeMLaQxH+XfxqALvvZb5pxy6PV4y70OIhZpZY3nyyTfVG6SvbTrmmIa1iQVX3
glp+Qrxenz5prQmzbADjjWEQi39nM4PGvTbdd8DiCn5on4/np+5j9KXH4YOH2yVhVk3Fo9z8QXrR
/iiF+UKVAhEZnbZLD4p4A46YX8Lva+zBkJhInwZjCbBnGbmv1AC7qDCtJdUfSE4rytk8DnbG7D80
9SB2Ny9/4UHxKRXoe6EObefI+QJz7cu/t8MijHtHrd7YLpWft9QOGZPRcHaA3Them6Giwvho+a5t
64dnjDaxAFpJEbM5hX3IZK/nmsYGp+oEvkAwcZyEhzN7Q/RYTzzYyEmn3gUE0Ph23HV8wDvY8izL
pOVdGukxNsZuq5oS7leVP1iEefhWvcRdcSiUV5ePgeCxgCw1zt0g8XqGp8AqYVYuNlPlbX3W0VGi
U//UqZVF5CuaOjN3qo/VtC+t1WzzDOEzOkkCvP9/576KY0mfxg4ywsjLEZfFFAhRoa6qSnZbMbmJ
rD1oMGaiMDrmrevvVP79AaOc//jqmCXTNGkKthsOE5IfroL24wXI5xg7bEHDYsHMZzVDqNngVzgJ
cqtZzAKwIVgTSkbNMROiL91OcV5GrA7qjasFOK1k7R00ol3haalsoY1bBCqtEVmAtUHY4IGOtHIG
V+V3sISSX26wHPm7JevO6dbMAvTlRyxy8jorYUbsGKHw4fy/PDWsdnF0mjqo7ySE8Ah7D5ybkfeq
TW9kwyiJ99wwC6MjD43ZjZVV5/9IH31H7TvNM4rmxuZ24rP5NCMTRmU6/8P2X9E53sVcjBKlw4o/
feFBVkwjELWa6LuVuPVO9CpzOOCNC5XcGRNxODpT15TM1oVRauqHczRqbcfbeQ2LlxC1toeqjoEX
zMbM4aV4EaxFENjY7yQJa2EADltIQKYo7DbjOGahWhxJj/s1EJGyYAz/jty8vbLF20O5issk0iJg
8QihIO15Evi2Ib6pOfuT8atO3lqZSpfIGnoGehgJgRJh6yU06RFwQFTjww9ZMyvAZ+b5vbQmztPD
TABGW7kfy9yPXXn0NMSuoeVUfSh9/n1HZ3ysZAvv2HymTZTM4HTOTPdW5uHxmi2YKPWudNr5lUXW
mVtMtDRHs++GNlLbshA01DfO5uM6cXfyqyg71jyxxpCMfAMcFl3x2inbX2qXV0wzPfrzQ0Owdklq
VZZPqgw625llaT12bppdy/5nf6RM87MPY+C56vAhgVHGCm2eCdEy8+UkS/0Rdqw2JOk+L6igzehq
wVB95S/NBoJ5jAJmkL52johLQy3vexlyOfFalTX/+l8iWKEGzT7rz+VgaaXhlZlO522L3YFeZk4e
T6GiU3jwSpFKIzomTXuGai9bRxvE0dm4idvbCy2cdhv9+/wutQBX1cF/wcTwHGdrU+eC9T2LVwIG
hvOQW2rfE6JeP/270a6zzqBpBXJkx/DAtfjYOKflUNVP8r3MvVPpCE36DJtp6hr3rV7VfzyXr7Uq
pMelUVNShYS8oPVgysX/RsIbOestkgU69lh7RII31ps+U2aPUweYYVXECL6xjidYtjARvirFAq+k
WTsii3cvwdXG/ouapz5I6XwxWG2LQIxadomw5WMRn6yUMBU3iALnlZUGttCWPCjTZgaSKsmCfmIF
KbCAbV37sQVSnK6hLAQqAApb2+kNr2/x0CUA0y3kqcEj29vAa6vglt+pSfxBIke767ZHFg3SJO+z
x/lR6qKCsO+5uddNsiYF3l2ynahCIUSJ34xo4ZTRFKxuo0MLgpPagndflOE2uiUYG9LCXy/7Ial0
qylvJlJm6bOjYGmWsHqAgok9RgkpPJGVQPk+zs4DVIzG8H7lB2+6O4T2Vxi3qiKEouXvIu+ch0Pv
fKN4G4yG0qZW0jugz/FsPAzXx7hEx1Wr9evQGAPXkBAvCCnKAV+tthpztFP3VVSGm+WK5j51Zzcq
ZqHJ5ssEgLS7Ys4vBTnVRYKeTzTqUaanqqhID7cHnQUSmI60G7Efhyvs7uJDf7VALl5uoW6NngNh
wuhQcIVHU8F20wTvqGWv4MlgE2laafgwF0pdEOEVrpVs7Hc1j3hXUwBMjuecQoarQYGM7KEK32Gk
+5DMM5OG4CA5VXa9Civ8kJmIbvs7bwXMyW+2LpivpeD2N6r6OQ0WluYiqN3uqR/Xo4x4QL8jtR0+
dX7CN9KQRwjY5befYY5L1n9XE/17uLgAThpdqIhzohJZOJ1L/nxQB3Ygc4/40Y1GTQyH+YkoOY0F
fHHMlPOg8xL79326DwZVzCHlB2WMpnwmB+MXpeeztMzF/RI9dhRL697FX0imSujemIvL7BkXRXxJ
MR2lkEMQykjKbW6ITcTrPkim22aNzTJEIFYvWmheRBcSBjvteNd7fsRNVDO+hya2AGQYfFVTLunA
1XZlC9mIl8Yew5VlzdFdOm+fUID/JyrQkUAhheaJUdgHELtG6kobEShA6cjbrUW+6E+u89NjHvCA
tGOynUP8RrVsc/dggrdtSo2fMhTaTmZwnq+CsF6cNQT2L92wj+rWsinMvnUC8XeMv/6gMTbWvtyy
Zq8YAm9KzXgXpTMYop5XZwRBu9xqbVzEOGz5Ct3brrE9Hi8KjlA2GEqdSwXK9tQkczk5ZYS4MNVb
1GDRrlfktS7CNuW6JHEXvH3SxGoRZtLtZs7JZv7JoiI6OX2IYD89315TXqbnMoE4Cm1NHPh1oSrV
hVz8JSR9v+2q1CvTU7/X0OdS1CehJxhPGX97n2n6oWwdVatNJoOM0ZdB3IDMy4flLNIONZkrqD08
1+TxMVtCxrSgF5RqedoTzww7rtEd6AEKNKHaEOCi44vrl8Mxc9C6w5ev22AWP+rejN5KOHhFLTOQ
3ykzMVlNhem4U3/y2Y5WeWIsUFy1Dq8Mj2kglnJadCFPTe1tR5jH9gIzqBU78ubpb78jVx6wfHX3
nsAbSJvIoZT5xjtp7QcUq36pz0V8NV3P9zWMHYlJ/rHnCbxGPyb2BLLZN8IhqDFmbC3mjJSL+wjY
/029NlkzXZM2wz/YEm/7PknAt1SAnWBwgo/i291KjNKT02ZOJmuW4eLDiFVuHhdjAnyzQp6/GdAt
b0SuKyxblF9I5eGJbNTs7DtLIlVplCBOnshKcf2w5d0z+CD38tmYyAYGj1bxBdHYXHdczPFLN97h
SnCOjXU4x/2a5v4DRTcnjYkfNHc8ALE64r1uDWiynnQ6mHS+8ZvwEDwCm6mbVxmOtPMhCr4uJ4ot
2L8R4nNQkPN0vXSqrVDKgpdW1hkWMoBgTUrZtzVyghacI88pKfhLleQXgs4rRGGP0+hJ/s5G4qY9
r0+C5iUk11Wxh+aoLbY+8msY+eSEgpCg/eXelj3OLmaCt+/Co8mh0vTXpivgshlHGRhz/oXiZ2qj
HxnMXISo86oXtC65zaY9uVAVehBlbxZoTdHM8zfqN4+01naEDBjrL+Whp5CZ1qNPh3ScltM0bV0v
9FvmSNlqAtDqYfxs0/fMQKHGUQu8bUb+jQnTtvaAM+5JnAnA0Y60ARtaAD9E1vdL2Ozq/hxHtcC1
Ap+Li67tTF6R4cA8zNuhTGzQef4a0AclbEskx3oiRdmhs3/P7pxIF1/Lkz6zJf0NeSgwWy+KZgKY
7Rrd2WtCH9yCLuMMEFh6BUQuX+ZbfQv+CCLnXgJBSil2bXTmscFP1d5ltm4LokR8t+TbGxuscZ00
WGVc5n0nwJ6CoILcr7GtXYLY29DoYYnVsCpnflh8kb3dPZl2p0SFuUdepHG1e6/rdeNBzkjH9xKC
91w87dmm68lFdPXOk4dJRZdTFJx5R8KYxyxjfYoMItWU96Ca1sWXWejmsJG4a6WkM0Pbo+G9cgGL
STQaER+eX2xVpgbEaKnW/+3smc3zp3SGhQ6ixPLhYa66bedn4BmpzAcCDBCJIDVrIvEPub4VJocM
dk1+/HpWUfsKTiscUxH21WeMfoCXK2WZTN8lIaHi8LxLlvi5Or6TpR1r/AmFiZ3AFusmGHYoXU2E
PzglaNJ2vZJYBtr6GVqsom7BxBn5Z4X2uH2cOJm+ztSDtlJ5P3kRVTSU8yAhI5JW5dGGtaHEf6Cj
qzP1uaRZAME1Boob09c8PU42MPQvxbUnHxx1mK0jNmerT3jS+F6OYgNVBELi8f8YKLgej305esQT
N3I0E5he4EIFnvvv0VJ0TpiitsGWc4NXMRRze7cj72JrdcWKQMCyJRlPj3LtrWb8n3uHIvKowK/B
EWCjqC/vcjev5Y09oi8dVHclhFZlPMeWnIme5BxGAKJU623hul8P+m2P3fHn5U+BlLWSL6SgW87O
afPddZ+VMYivYVMMlcPBt2RpwB2AYmo+YOeWxkMFklykEErvSgTNewXVF5niHED9SlK3SOhds8V/
vJ2TiFUnnOQAwXR9L2vB7+/QxHr7piH1tAO+Zj9TC+0meKh9Zl/sj5D2dJPFMWJfcaQ9dQzq7ZFk
iFQPEdjVUb03hdhx+Gn64Rg1sobGIyRkw0R3+9ocFsLiUX5rV6hfyvyeN6LkToE8nGX4tshiKtQU
QJq4hJs6SM6GT+TTpkofCz3/at7latc7vD5+PILUrW6Tq71jjJlpEx0nQECOjbCfbxh8STJOPX2a
Hc+hWt/iGa8ErtYhhHeKjhOPIJ4J2ZuTdFtc2fL2YsdfQjJPRpd3LimvosExmNFWZHJCzF1J1ICD
9Yv6uQhT7q9amm+9+g/dE9TrplElEURihWJgHkY2fuDO+r3IEwRBCFww5PcdwgUH+OcQyGk3+xvV
5US5PrXF57vLzeltG78rDkSDyCFBaWH1Bz8qp228Fc8pJT2qy3KYWyD5x9RVrXRGLVUJEfdUGR5h
7W1FwyqSllGDNHiZ22NGb0AOLRL4QCmAUQEP5xuJpFCC9PUHrPzvnJOV1XFIZOjQr+NvCq66KvOo
7J58Iz75Jlaaa9r9LMvAMvXjHZn1xT7j4l3R+h0Y2VRHC8OVKc2qHq0v7AaboLbPAjo4iVHjcIzU
CaS/HdlOqSnoUVMjW3ZaxvTkZ8fnsWf9Q9/6WWnEpIg2MzC/CbfviWeqmJordT17CckR/ZMDgq7z
fB0Q1CWUl1wR9BFLsk2GB7HHaGspJIIVzvo2c3WOS5iZCpcFQN4vXGUNvQTL77yWlyVL5rVOGAH0
KWZ+omQjWom+7uqUV2kmFsDNvqw+To5zgiiIj3edKnBr2FM4MBAlsqpBCPmO1EVsv2q8TwEiIEiq
LurndF7O3LmtLBVbjNw+1HkbsTLs1FoffD/VgLb1g543h2QPTrZLc/iPU9CXKY5peKwme7k0wKsb
zeGJmjPGjPYAyEmSyTEqHBysOf5798B93ZrIVoMVTFSH8c5OMr+GLq9b8tZ8DahBpbXPcU+0qxtk
mZM/suWGakISTs5DiuhED+DuAdUWJqCjSY/JlZTNGhZ7ep8jmdfL8x/RmH+TsA2VedE07ZgcwyY5
9Lc8kw9Cid559xVplbITalGPcWecLATnT6ApgU+wpQl3LuPHdjC6uAsGZtoD+2Vk2etYzu0O6HYJ
b3jbpJMZbA+k7CjMrJyOBuyj/P7N+sPlkiTysC+yH9Iz5mVLuy+VsWXN7Hl8IuS+bvIiuSNIZnnd
mATRTXLKe5S0ALw45oOflIqea5+CtxpD1fYezV/OAWMLOKlK1hJcH5pWZgq99FfWhZc8o5dsD89A
tti3ZlwqJaoVZT+G072671CHcywxxcfDF1TqPUtImzeiXB8+5AMkiejRIQSLnA75QADORD2yzb3J
3fQbz4fMmX9rVIjlj4TWfujPEJQaHQEEKzAu/gOO9uQSgQSCwZ4NxnRJ83Uk8FzOlLw7LIRTeg1G
K3bEBVZ9A8hxLG0HrHZg/SiYYMM5izcKPAhqctDfPnut36xPGbdK5+Z+bq5MQt8H6WBP4PKfDy3w
bBrOFZh+Hr7IXgZMqi8BFW72RCHWiLrpey0fCif7Yd+i7enOAftOhQ1vZLp3W6s5qEFAlvjTfMJB
KDmL9arMaGRcV9sBEc/CVgxdUzd/SsuZnmbbRkD2mZknQx+EInpsWnPL9V8LEJ3AjzC2h32Ajb3E
DVJeoUiDDd8VQg/Kxem84mfM3N4rhdAx5rQi0hT8B2mbY7SfynQlF8gRUZoSwm9QJ49m9OlF6Tj7
+dMKh1YUG0I72ykx8yK+yrVm0v7svUt/smq7GtL4KpSsvWkqVlkulH+FQlKeH90sjJOh6FjCn4v5
4roFbRodlr6dMtmfeGySknF+QoiHUX40ymQpPFqn0b2IDOhc+Ci1jemk6op8rFSQEbqwlhVTv3nO
x3LTpIfSfOmFQjOPUKUgJytg1v9xuGENXXqMwcrykd0tlNMRNu0CpQL70j22leRSAdserHhq2Fw+
DzVr3KDBjQF/8MZiHXwalLEebMuLBWrILzBxn2CLhAeFneHna61G8tDdarhfyP5rXp0HorvLjT6k
h9RfiJtFiUr9NiP/MG384bmOHHlWnxCCvfTlYY49A1H0y6R/ED2X2ON5piMV0XCLJ7lnDZ1hD+Ur
1UcWHHSiFKKr6GgXH9RPTKCr3PYdz2MJ+naKoUxRSh2ekOOIWUhofCNSD3yddBHyshN13KTr62ZK
UUr9WiMm7buMtHGBFKKIEc18F1e4Ja1hRT0+9ZfmFjwfhTSQ5a0rXCx4hudj+V4IKrPA0hGuhrtq
Zk6DUDuwpYwXe7jeFpLywpn5D+C1VrpzK1TwmlU/iOyVqBb+CPsjUuykGZnIALoCSEXg4Q3gJ0o+
yWag0zT897lA0Ex/7MTU3s3+SThfABfsxNvZ7bri6pPv3azNsgz06DdJe4VrBe9mrbjAS7YvWuwD
oFNl0S5qW+1PCd4fmS1+tKUc42iNoD7O6Q9t2Jj3enngY4ZKc40ZhBTigUFfn+Mimuc2bHUTu4v9
5s+P2VaFZL2O2qHY6xXYoEPPYrCw2/Hj7Hf7ffRkAnDGMhIhdvu1Qi0mytBkdBbFGftuRovXMOjB
1VMxRweuOsLKcJib9+Uejfg3R7FABm2lzEa3cKHAxmw1VLb9TbFYLQSVRP23tJJ+0/KpbqVwihYj
mMHDjUfrdm9xFtaRjauAUXKgja8lp4j5gj6I1PARvgzTSTPKYrG94urVnPNN9dG964Nysk/8k5mQ
ylOHAwbLQE8q9ySZm7MtoQ3Yz7DNhjUEQ3rF83vCmzBHM2mSPQ3IC8ajgI++2C71ZFJoWDW5leRb
An2E3C4LsMV/EzekdGdgT90XnW3g5UyhFM70L4ItaVgCxgSUAX2d5dtPnw1+W/2kzdApgjm/I+yU
ducNMCflF0nKa0VAQ3N0wX49avn//5EUymLqGg5Uk9Iewapvcs1mIDl20peysSol+0WIt2hn8a6n
kPLzRd44+q+bYqOxZE3W6YEy3QyuEub/OhYNmBMRphk0LuBYE08z4CGAgEXeF5wkX6i/4jFI84W6
3MdviF3IJW6yKtxrpA9wpEng1JSMTlwRSfws4Ky2BdEI+Tzfpz5xomeF2B0/hGZ8jTidBN/L1QMy
b7L6b2DCx3GDrFSqzyXpVjRY6toPjKvLUxf/c3Dq2xb+2tCjWQLUQXoK7Cxsc/Jom96h7mYbJBXd
IaRVg3bNGUbcMpbI2ZvjzorlPfnlo1UgSBg+gYuTMoVe7XDu7htCGLrNoojo5sx6euWuaqZ7m92M
dCJ2Uhx4R6GmHCpljCzoYF32It4h3mbcMIZ2+x6yEVmI+cvKFLhqfF2J6W8fNIkrzz4sf11OkxXP
EoNdXK6OgY761xPW8SlqWhw7dm3NYKGxuCv4dHqWddc9RK2mD+/qbBj0glx1hUZ/Vt263ZC8HVxI
XlN5JcLZ0zwrqwVz3HSUvvmEXFuVyp2sUNaZbCGFi0r3sNb+U+aHkGSsTcNl+QENMZqiF+JYrYQd
gPLoN9Ipe4EirkWxl8mXR2RNb5HRRTwfEdZRGCRWUDvZhlnbPIlxra6fXepT8Dr6ZZbwArYX1nwV
z74FrkgqIuGwUEZUNCP7fhzrX7x8KTebO+EINI6coiwG18HvogZsMThIhHAP9Dq2q/+pwpvI8zC5
d4mvW0z67rvdhwtnlmhyLrYtavxDitsfgwBnElNadm0db9PK1d+v4vzIi+uzfZzA7+/xFzlsMHBC
8Nbk5e5rLOgeLHnH8+uECTCRHTvQS0MJIAS5qJwCdVbeOj2bWgiq1dHet/mZgImLW/XxmImw5o8R
fHN3wmc66E2NBdDiM3YaOxLotG2OZPPDCo4qMTvF80fnywn3o5KjROgmr+wr1eJnW7Xo5jimV7gu
GjSM0VjmYjTRutpBcNWdC6i5V/V7h5MASQaLqLI0tb9pnBOP2/22aXarAZWtTdhfrKlk2NDXAe4F
giCpa4AZuofrVCkwRA2cSLhiWPiraj2StvC2ylOFdTTTFa0b7pUbfFMUFaMe2j/tx6P6PN93cb7D
bSLY/ZlVKkC/jkAWD92AkholSwmJ2v42nMnnbaWRZcxfJcylRm6TVsG6/ExgrcD6+WktMyKuuRx0
6LWm/Zf3p+UO0P2HWO7CXX5dZrcHTgHMWkQu3YexX9TwCqpj+Jth06L0WJfKuaiMlFquy9yk9ul2
NJHW8bPz/9cmMogIJq4qkcdH7AztMEERlcTd+R7TSVjK/cIWLBL3qNgfOIIJcFVb4mWXh6shJjQA
1VqvUdFwmauLFbXeIIjVx9C6yJb7WdlCyVhm8ibZ2MXOmezSfq4YcwAPYwsThjoF8c/eUx57TQ9z
kbOlWzdOAkuNFGWIoA/vhKwjKsKJl7BZb48o7Rh6Ru5HgcwrUYRZ3S2XJgiAptFK3AJPuBUNP+u4
vZVd+LulvEr+soo6PoDnz6KGBsYelOx2d/sPFl9gfWYNOMM7v1jwcWnUFR/Q/FQOPub8QMuc9zBd
38wmJLPDFSlZse537kO0UD9jl+bqYXDLMV1Scof7JbufDY8RT/GwesvDJR0qm9BUBmXfNi/hp0uN
//WWf+LF/rBoyeHu4xZYw0AhNFryiHzTgtK4ZJhRWqc57842euOiWs4jKM+AXzKO8i6jT+9gMT/5
Ws/nhujgmYXj+w6UcpLlfwMbuic1VW7iQ9wRDG/rsnoK6q62GaORi6dZo4yUssqljxJodMyDdFHX
+Oi/m/QO2jcHXEgK7qjS+Pq0BNWg2htqUcSp8SFWKOu4X5JQb/fyeJw8qzPoCKvTGhZTgMwq4hBf
npzcTa0gYj4E6uRfOLldSpmRq6RNsyl9liJ7FcNFB2kztg8C+ALO+WJuNojBzWr51xD3X3tqKjwv
il0FTmwfo6fD9mBRWg2gdAQVDhb+i6BkBwu7GswwILWTA6HW4jY7Ys97xJZ5klKOKRYnJvJ2zwge
gIYOxiMeTVPrNOq+n420DVaKYz20ICS52p0b6UWJpQoKFeU53Lf0hlGIwPLcZKuW3CSbYHU0VN41
t8XdWNgKEekLrFwoPYigCBWF/V9cu3+4QCgFSoAU7XP8sYMnJY2agXV+W84PACHhAaK6naFTFfeL
KI2rUlOxSzllxbWp0CQePnMhk4Hh0Grsw2fKqDDaCmxlKsZEF5OcaGBQ076CkwcUdmBkUQgSlvZt
6xRbet584h4Z470OmbT/0bBqpG2VeH3beVnRdI1MvHucryrhiGz0jEy/dgtB5BTDM6Ao7rTm9A/M
x4BwRW4GOQCBmg/7U6CneGLd1S9dmIy8Z009IkQVHKuAex/rlKlvrx/Wy0+fJBoR5OZ5YhhwT0eY
MbW9ZqzgKGc8SfQHk21oiw54zI7+TZD4QDNOFyZGAzK1ln7pdBTtGu3nqMGbTY5i8rxlwaRH94vw
uPAGoWVmU65ZNG/9qG7WhmqAbJ63GapjLyqfm2jZv0poTO/U6H0BQW9jF0k9LQufGoFCvsZE9VpO
FSz0AC+YaixsmVDIxWWkwRCpMHzILcAhLMtTAuJ9gHz6Kj63+u/Ye0/FJIVmNIcXafA2SY5E/6Zv
EJjNcpp02ynenMn68bWJd8TngM9sieAh91+tDhTO5gEq6Fp7VA82udix9+zNz6PYd5jqqWsDO/WS
hoSnDcF7xmNIifvY7OLwPhSPO1fbhcYPdLhXalNzTZb/yw2thdZx8Xr5WqjoNnCMhQqbToZwR71f
dcYs9ZBw3lT9IWCcyaAS7pBk9dPIB7UpDHUoCL9QJooYjNzcxRuQljAq2M1S/kbtAHjVqi4VHvmQ
moocWaUDiy0ZDDpgOYj0viX91VtOPtag9Szklikq+PsILlxq307hdmlboUQk7SwW7RXL3s9oAbc9
nDhMPZXm5mzENfqfPVQdA+Tmb+EDSkAG9/KfCl7BJB4hfRf748nx3sib9ubEL/QiXAtFofjbJBgu
hzonTEzfdBapP4mwyW9/Nzi5oKF8oA2WcBP9xN6kyK0q6YDPVt8McPEoPrw2QoNMMl9k8vC7/On4
BqfLKePMHltHrCX+wV3F0dv0DusYpbXdxv6aT/lLnqm9eHaigGqDzfklYkmhGSjC38Ad2cAUVRZc
x1WgLDEt4LB/m69XSBKVdt9I/Gksd90nk4tMNBv1rYq4cKLpMhNL4xbAOwH53HVnzpvTP67jY4He
VjeTWGbsV3cvuK1eJMTj2hpG6z7aJuEWvv+CXKQuW2GZ7mat8rD/lyMoHlgZXzzh06vembHaFcRf
8PBDs4F2dQDoB4If1rWtUXvPZq9LjAWOUzqYs3saWgF31dNJhy+LeQTo3sJql2Zi9nX0QOTVna8N
VNsziBvV4UPlGnpeKG4D3von1pgb7tijJI/yT6lBYUJBg3eNYAQ4P5/yjrqyC+BB8U5ejXwutyZ2
CV2dUFv/+FVHHS9pnLaMM+wCmPjLHa2lamm231zNepXBPikyUUDvPwmv7AWB4EZ0zC1Kv53c8+/U
OtV9Q5ikSyxPVWhTvMAlSHcn+xVyl+3tXmmgEdeQ60ZxEE1iu4x1qZEaQUCy3PVKO+9IKbQG11x0
eFBTp1i25DPQ7Hgqpg7cJXHCZ6lqEEvYD6/PcQFMIRl2orKD6Vqr6ijSke3MqJaTO3sWK3q1D2En
HVL5xJ4ykT/XbreUDuKjql60NknSwE/st+HncsN1w+eM7F0fRsTCdwTrWkR2mXRnvDYd33w+AHUX
9/zfvdGhgZAh3H2P9874lPQzj6/mxi4rCH56lU88TlOaROJ/Hs3Np06ubpMWtU/f9nC2qN9XyxJq
T8K+yvEFNYji9V8r7qjWPZlX2HGghlQa7AhZO9S7zn/pKt8wwGQUFiFoaZGBtXGkHNfWq1QNHfqU
3A0AJoEOn9WCs+aPqNLYUKWtp/IiPwFh3Owa7KHHBiTEekxqPZhXwpFeEb8isZisOrYrB5xr5Ov8
a9D+aWlWo6Lmf+SfqzacPaC+8ibDopXN5lX6/K21qB0LWtVoeL/y/x3Z7NmDpV/DvP5YXBqwqlqD
TPvZ3L5ez4HXjTeFBi1HQMs4XFLEqa1dR+6fBje+oQBTq6igs3LeIG6QBPymroJ9wr0bcEkRplN4
Sw40tiwkkK2QlxfRGegWbz+A2UaCYHmDqHjOaqiqyYopNl1kUJQ0LJdqvnyaSfmyjC38sf5iag9W
7Pix8YaJKAWXZFZ40mXyus/HoTiRT+ko/uWKd6ke4SLlPDx70BM0MHSyiro8kO2BHTtn1bPQCg2a
u8uyhbFk7Z5eK+oTPtutnn8SfOH9LKo4Pak0bUntPAZ+vt46cVELDSLOUJBopNF/NqOhnfLg2XlZ
qfnpKkFlxWRRB+q5dZ/gXPJooaaOlQs6dMlUByHpDmfMsYq5yQyw4TO0iTX0cd8oVTuFQ+HfJxFN
LLQPTqx6CEwEaWsPct+MM1Wt5c5JWMG08d6eRspXwzaaOjAImpekZUj8ovtKTGtCM43cKuVUsCe0
9XqIb4SZY4Xgt6bj5naXwa50z6PoyePiyVQd4PzTzMhrQV02lJmSFW1B8FLqIJMAOv0HHW6ltbRS
3Y3gMjO1qXOck3XIltAVMLsxadZjWrjeuGhHDlpRNwzEht9Qix4ZdP9LbiroNt6EHB6LGxPh5ghQ
NYhn7yhvL8GraShWHvIRblKJvCiODFtG04gWTyYVrbAEzFOOGKaH7VjRWPEazIXqXWsRi+TMqAMd
vKWT7r/9nyt7K707xFDvv8EyLnqnKvsDufk8tmf1x4LvAolDvmi/+YdzxxEnjouQnk5VvHhmTKEM
DZT95oM1tLPYoqD+Nsw5PRcrCVK0zPteohTbWbkQqzEoSlgPbzF0b2TDg5OqCJq886UdkWa2u0bu
onK4p8KRQh4RbHBGc9VKxj4wEPr0htc5D3XrMj182CjHpgVnrJoq9XwjnXqsRwbRwCtQNtG7qWcd
zWlWeLsft09ZhV4RAUDPoapt4HGCRorXiC/EUel1Y37nhiLejfuyEa1zVmxvAYNC98oTRoUE7rgY
moYh2jZUMxZuXu5SY9OLKUBY5L9GM9D9uVl27g5DrIFmqOI1ZCqZXkuKfgeC/9T9SXSCIvUBD4eu
+W84/J4iE2bamPvHUvrh2NzkjTdHrqRCoyHc+KcTQ7kkTmaH1r1ZgIIRWiDce2q8Of48lBttMGDK
cdf/xpV2Xzk4uzYG5TbeMDSGnFbIfWMqjdHAVmmOMnLxCrFWmyC2X3WwaCTFB7XZBn7GNghXES/y
XTqdBF/EvdOA14FswnbkkGh0jVECKMlVntOKY2IvCAOhiRxOc3d1n1QdjBS5mJQ31C/OqiDJeCLV
QgBysBz+nr7HuNFfpjDeO2eT18iJSctt6raabebup1xxiGdcv/Om+soPARRUsdnhbiSUFcuC1plk
ZEPgzbSeVdi48BUxDQWrFLWVxaMFLqEeTrz40g6OSxOxC8uBPrNnG6Gj/ZDe4p0SmkqiCF7hEmOe
r+8Es5vrZ6nisVwT1qpEX4xPxibWqxrDh7pJ+wW8WjO1llZOn8TceNKCiYmhTFkxq0CRcJnZ1sEA
omCO1qPSLW5/ybJaphYh7fmcgr788JHQnepTP2Wu6TTK6dNIkBV/fB52vFfX4C8sblQ+5utU5RvC
8EsdE+Lxdh5pjgfPGWyGBTjPoZN8gRJtte6qSn9sYirhpa2ZrgxutLJRWs0k0Rx//mgR16qPyYGb
9NAwEKgyX4/Gz3eAlzA3Y7WW5BA6AKa72AC0uUVraLq7j/g+tara/RQAyEsp88ZnqyU5Thfgb3xm
2Y+uu9wIWZ2u3Yw4bo20goDsWlLzB1cg6njAeNxTZCnW6Odw1MpGUr2D+gWzx7t90cYCJ2AfmTCS
7gh/Y+qFxTFLvAvmUpouGJcSP3oNeyGngMoCzwtbOLbkhtkt+PGNVGyVWZKRiZjNlBkpIYXJn81P
Ot5qHXorKb2ms9aoy7mI8PyG2m101mfI9FEEYzTqYXl+pr6DXSzDDaASceR84EGE7Cx3TJY7+0jU
WYm2OLnsIX6H1+WgxyZJQ4YYxYpt2kmroQctheiRCN5+19IW3t+yA0VIF5uoNYDXv9ExuuIF0eiV
2aTdpp0FWJkEe5LWraJV4i7RDNK6O2+ka9ne1AtI3haXu4oS8UPQI2qtyTkaIoy2BjA3p1kHGinj
xn3Bo7iVHdANKQIxmLdd1xwCNhiYe4Zs801c8hZZ9hxAVT3vT89WZeNs+kctTlnKUxXoBM912IJD
S0doux4/+h4SFQiuObD77h98hD4Hp0zaVkae4I7S9kuO6oX6XjBVLkvwXj6JD+mfG7mzlDfM1a9T
HAlMVs7DD7BHX03U6QNWY8Go2CymQgQFRxZ1IfWVckqgrOxarDFtI/ZZM5uKu0NUpMyH+ZByFjUf
4a+2+71FB5r6I1Z/1HSK4twvowfQzTyXc4XcLM6mb07PxNCYdr9iud6UjWRoLQrQK4fucQEz/hrd
Ql8VsQRs5ivF9PALiqfx0wuFwaC2FkiJqNTGc9N42mf2Gu1IWJcCt78h+224htT8DUUQxXez/5aG
QvXm++m9iGLhlxEZ56ZNpgw7DImINlCbch+M0EyOy+j06uJSHKtzi0SVjJamjM19xbhK/fGznghX
R58ciVYPI0SrC1eyHa1vQMwccqZtQhaXw2vB9wBAhn+qTNTMBA7DJ78CspYBb+pIKuYohWntKUK8
U1D0K97eaP7aRykit3ePSLtZMj6Mk2k4kO/3FBxbhDn9BDfmuLyf4vyA2KFA4T8Yu5s+niJlYrxo
Nqkk6+GXqOtQewTb4MFvg5Av9uAhuNSPliltGbYqJuMIWNPcv9Q+OIMwPh5YFpr0ohrnjlUiFuOG
LTpD/b7baGqarcAgfNv+1+AksTkIr8PjpcwWjBhvy/gGX9xuLbRdRLL7gqWDcPDh18VIXuSEL/P8
Ktc3JHts9rJ2sZn7ZCjNz8325c+wQCqyngKrqr9K+9/TldauSlWNWi1ZRAT1IuGQdq6BykSs0lFT
+BN89V/Wh4WyGmVXxLIc6/Fu8fplUY9ixkn61G3dyq/bCaQQEnrJUhsnJ2j7rhXFBmIu3G8gzXVr
uDdremMSz2amN6cI9E6ZhtISnOHX/ZwfptzRtimvKjl5qE7DczvUEDc9aVhbZOmRKdPUkV3dizup
+3I7DOvvTOO0FepXIUNt/+Sj366wafN5ei5ilyJ5H4VyLOQ5JqbAZ0jjm3XXEzPe+q6NhOeECY0T
wqPEQQz2uvoumtYlcsbg5i6AHHCCzDFVIqvGulFxTblIkRIsZiBpDxQ33Db7Yfzpxi02Nh+bG8d9
T5xikElmOJ86FTiznCYrnHOtIuCV4TlH+2eJxbkc7qZ+aauk6oYy71tpbw+EY8qpuvO0P+5CIE/o
HHE+0m1fY841WtHZYM5inR9BSQXELIgdJm04rBDEDmGwr5cvcRtv/clshknvaAlhE4lnBsO2y+7l
/wCUw5Ql1bWFCK1VWrF3J2Z8x8QSidJ9DxJoGw8NP7ljGZKOnFAX6sbiHlrnWjZ0Lv1BmIJOlbh+
pNjSifdAaR+nJlojmvSuAfx+NCBDDn5p/t1MCDnTDT86bKfIfnjpoFGCtSX/AmEmqAEnoaIlRp+0
p7PBijcjzryM9DR7l7YuOD8H3I2nWvbw/Nr1BVuImOV7dqpTGHL+AVRHyW0saqvCAwcmx+bxpgl6
O+i0FFPnrqPykzUyyOXCWLX3ihAw56d7IEHy/nZwIp2YzT7W9u8EVA3pDxvr5Vzb0OrPMiB0Mzy2
JLW/om331V5DZ71Ul44lJok10ROqIeHuF+VZy7vckiaTl5Xq+QvIabfDaD7FsUzXBtnaE0WhxcEb
YhrQMlmUTnvoNWlpzxrZevLM3NsG+ZDoLSBJmJN24zaSlZEjkGEjY3CY7BPGaD0ArAQ0Evl0nQPl
zJC+6+qmeHflpyfcsZEeIZ6g0TRF2GN++QFshbC7GmSy3Y09vFedZtKj/0fe4BHUSSQOxZZXMqM4
NG5tpSZSVpR0lQnGFLVhaR8Oousbm9Ko+jCW8wB8QhHzJqNIfELNVQ9ZjdjreXMgumCt0zG2dPyV
GcoBbmSC4YaoSA8SgW3K/0mv9sA8QviD0KXppDtmbW8tXGkpIOLlFj0JojHsqs//rmSMxY5y60Qq
uNKE62CFYDgzal35UbDTYIXg52Ydm3UYaIHOWS+rAqbu0zc3qxUqQJT/k1DwVm5XPj8NrbwfSOSv
LBDK7PhHaizgQWNBiLFgMTR43PiiVHVLbnPH8nItXgR+GbUqUHP7p6vSS+4zy3JfAZKvwoCwmZK0
mDWZ3w2cK/oJBehL67HvNivmT3yS2XSYenVEmnldhDElhK5tDgOorB7JYPxVZOqBpYmO1koGszJ7
L5ovz9S+Y567mI1VNf024yxhzne0cNANlnyqIZRB8uZhPUDXB5vpoXJ6oduzPEHrU6Y0PZOHW6hC
Qpf9S+L5pWeqwwcdrpMRnFcJDFswxr9J/3dDXklnkDA3fQApTHC72Z/+B2Uv8Eu7j2TUScQp7d5U
Ekqv1SVf3RVPZrXOOnGXp1VyRsNCYnpf9cgmSJcd7gQUQmVgYsC90d7ywyeS7l1xy6SNthJmMMOC
5t4JxjZiUeDypkTy58wRx2nzeSHAAz2x3PA21NruDcqkr5pDpzn5lZIjlAnEsI/fEoOD7CMkGvLD
7FBN7xvPPlxGN5+ZrF6T/hbQ+Dbpif3zT3eMK2+7PIM+83kTLBQALzzH1xSfmU8bpSmwTWNZMcHL
cmllF6txPYbfGftZQJWOzwSUqNZfHpIX7q/UED8VWVNszYMyxZQmYWyss42LAk2vOh9F2ontb/qD
YtKOb4s712qPHtK+0FTAT4XcH1/ZwzqvxADG5UgL25mcDHb9IXXJa6poT9zDi90FF8AeclSV9q+h
NyCjZij/g6GBmGGK8/L4xrGiC/Kn0Iie7qSthM902TzTK00WLLcIBu/Av9PxCceLVfh2fA3mXdze
jmwtd75d20e4vbi7uHNNX4uUp1fgPcLV6r76rzSH3Yg4kG91YGQ4l/ywcNc5Fp+gu5i685fQSW6F
7r5pl68Lp4cwGc2EmFaHUOr/IIYH6ODG0OlqozhJMefgs3nURwLM3DAjW8jOQr97izfhS8issIeH
4ymN84EWAmn4C0n6IJb/CL0va05IHcoMlOV3nAzZLox6GGwPyAkv3X7Zv6U8m828qNVjRbN/3R+X
sDlrGt03nT5ZX+1RitCwPLS+wToWwMu0iBqIyw8jF3DlHNlLDZHeki8pr/cV7YjSnLzhERc597Jf
e0W1xixNRqY/wL0QFbc6M9sQQbnlBxdJkpF7kC8COqsklQGgBHppiN2E4ZO5xI9BZkJGy00Ap+XT
gmgXyNwZsCKRTKpdD+urpOIw9niUSSPolPLic4MOqvPTGPk7zyaz8BEf5onQc8cblsn/9npBDcSd
JfAyi2ioLwhiQ71ZgJflWj87gn4+gnZnR3d5WmdfrYrKs5jnNP78p8g/73aROlmuEYxBs72n9wWF
aRsGfA1v4UnzkinTwO3mxM8FfPIqAEGgEV9oyLuRvqM8CKixZ1Xl4Kn188s5Tb05yOSfc0yxUr25
CHRJnCSVdwy53j9Ir4ftIvBD4ZruPbVUx8WVnq+qAL8GyjRS0ubAfcQTVBgDyRaE5THkpDumpNdD
nFqjOLJfx1vomymB4dky4u6p9MPHfJyNg4bufCccKmG8XM0pEfgEV5X34tZYMbEpiN1oAVD6j2H1
yihQjJkbGmTfhZvVITlyFMBC+K8JwJLXqjmQlg6i84RwM1nq1f8QUL4LuQxmSKWvzjyj1fES1SQG
KK9HjV/Tb9T30ANra5bgaStygF+Pak5sg2wm8Um6oU7qf6u+rBe6DyFJOeKnRTjkZJ2fADuLIXe8
MiXiMZum7GB7ektAzRVV3hLVjj7EXdOQi5twM5Vyl/QiysExFJ+He9zsrMR/XYb8QR2N5U3gU/qo
8bTLw+pMXpqgfM1+Xg4j1U9SvvHre0TFvbwZqEifd8sXF7RJM+3bNdOudqCcxaBeKz3HaeQhfGIc
nL0d9k3SOCtchusTpK5WxJi1qJUuW4qBGRJCPEX0a7HUzGL5B2BNbAnrBkjxlnbSKWnE959YWt33
MrWktCJLt+PtZUQm6RmgsbrpLfVcSzzK33aa7s2IbjSZ50/ECRmBdqJaLzsrAn0X0/XoIa6QKVAx
DKjEW3po0u2MqtPDiIN80UchC92QbxVrlo3ibZzIq1II4a5Poh/R7+2rKxCaZ8vvv6EAwr2nENKo
9Z32d1I+z3VRDQZtS6VwKI4JzPQy7KScS1ia46gjxUjWoO+BH1JCYmrt4E7SnQc3XloaX8Odiwkq
8BJVaFd+xounFBIEswerclwbwSej5/qSz7g3jK4smzncdKrdP795gZO1cQZwbhjlajzUeFzo/PxT
e5vZWmRhtEPX12sTCycsmLsLR6qOtFsgjDVv3WjZRotcFoHQ6WuF6aYzdtq5Y3pg3FtfM/S3LtXQ
d1Lk/GXu5oIhQ27zgO9/RD4yUq5QceqE7AsPmE+03t8mVl2/Ghly8f4EdfQX200SrQ6ZNCfXV+Fw
1+y9yujx0Mx8al8WmDWEdNBkZrqcQdUOxZ0/NKmuU6I7KeBSLe+gcC6On4CJi8xQEyT/tPPVD8uG
UBcdmgwh442NEv6J+q0zlVHrEARQcIVZeh9Efizb+Lr5XKBdUcz41DICQtX3Tkwiur+UVYGxgD6g
OCg5R8sui5Ow5LvLlbUf6qSZfbOiZb1qGzVS4OXfe/7Tn8pweIaI2tCXc7sgC7skx1sp6cf8/IO8
g2JtQQv58s4YrSqRQheruFVJZRorl4EgF++KuxTr8FB28Ae+qJiPMw0f5zwCtuCN3JLlu+oMoe2L
dEBNmzVf8JKwi5R8rrUiwQmOaO72aBHV948+2uNU9RWR7qSaXJJUlaXcNNu49s1ZGkGWiAQeLonw
svJCQxMojmtn79Hz/Ec2zFTxgcBbDtXlXkaTTXi6QVAv88I+wOHhOojwhOJ5w4ncGxnmSDAVjpGA
srLM0tlwr6sF9rqdL6jzYAT8tdtSHDcjp5m1r8v8CUW+fwvDPIBsepRgBwH8r9KxRyYBCJshPwS4
U3kpn2KcRv1Vz5kGFg+M35IDsJNI+eL6nP7HgUmQTmIdp8oHsGAw2g6X3zEKwIvuDnpHeKE+x/hf
SR8M87RSDahBB9VT+7jEsk3gcoR4WrhCNvPIxR1ulRLewo+TiQ3mVSA4NqwcNoarOsHP2oILVT/M
Y8M+dZiTHswojtXqnoSH3xUpsfXPqTVkHOGDy0LsCkTskhyku43pdRaEoLVzyxtknvWxKqBDCk6w
/02qhRdv+mPU8l898MpmKLJppTSEeI/MC8TvjZPrfv1ZmMfuVuWbaW6m8cQLz/g+7EtQ1c1FlCSh
vgyeiwMYnLC4jihNA+JkVq/bFfPHEhaNY0aSmcnHVUm6eF5+Ny0B0DbIJ4WWcE6H3+0f6l0wGy59
EE5oLEVQidivLBGysxI9mgy36AyZtvuM8flq1BuCZhim9cHW/IawEuxxDLDEWL5fqWRJUAbHE5nl
5SiGTG0vI7La57C7rjPF/GAJglAYEv3IajbA0ywZFeWTJbe5M4zT+QOXVIrGK+eih+0HccVlXV3a
kw/h3aeTyx4idOoJDloDVb4m46fJHNy0dMcmWCcwWCWYp9qYzu699d+nzXMhgWEKeYo+46RyimiQ
FV9FOLYi+2e4elO+podHWARNUrRqOaJQBN0lfYXH+NcL7kB61JiPj5dKFuzVR3LxJRvY0VSG7fbd
cRU9zs0Xh+eUiVby/HSaol88vj6dOTRuO2Y0nVB7DR+xXoN7piuVLxLGqfNW/iSn3uY6u39g4LFM
g+Lam3HK5nmSIQ+IXRzTuA/kvSJ5dN42siHMxYknGCkYu4bpHh3blxNK7Y31/vbOaMrQBMgEU+yO
s4bszudgRsjboOWTcs7tVKAFnRi3Q5481uyL3W9pdphgs9IOjc6oK23RjQXJFgaw65bdIdrvhRia
R68NhaLEO3ajXEsJmP/HexEjVCqpN3StdAqs8gG2bY30qF8UOLL7b6xJSUlIt+6Rl8woEN+khi5a
T+OVeV/o3Ikuyh2gAI+KwAxmKEfI5g3u0XY+SmHytA8GMmXOKV6BmHYovUhWrV/sH+CKgKhZctxf
Rrjd7Vglo6fQdDd6E0vvtQA109cQvlrW1TO6+Ck1wfMbEUDZAH+MbM5gDliwsRaNYwoHuK7CStFM
6JcXpvDankfxYYB6WfWGVS9lD5woV9vfCNWCPQxZKLP7bqgefZAWOgVO8kAaxcow0n4MALU+vAk3
9/1VyHuW8mZ13w6ftA+GnHdfSw8J7a6+i4S6hccpEnOxU8DOcqn3HUdcNk9R6TJYmLbRgobTCCg2
USB+gonX+gWnykCvJ6hIpHGEyrm2Av4E0X540yVC51DnP73zwt7Arnrw+JinnDgukX9Iv4zr0qUm
3N0Bl9fWAlIy/Zydb8iLLPikD4B57HMNhY3mstHxBoB1eT9AOGc+mt9/3EQPNwnio0qMn4HI4KSd
kpqv4OolNkUCeBSwRoFCL/wy5hb8N3xKDI+EZaVQClgprJ3D9/3IJ85gWpT82mx2rWpMcsZhW7oC
sjSd8HdNJEQ6I5/qwkGTiO9sriLVDdXAVyjWff+/Isjm9xX2jQCV+y8r0S5sQxxEhAVO7YB6zELe
cNdWWBnDweAY5tgCNaouaW6ZfwtOFXPlxEwAL/aTIIy5QF29da9+unApOm/dR5rCtW8ADMh4Md2e
qFF2U96qwetY8fUC8S4F3A9LzzBsd5nJuggmC18NP+CN1B9GwVEedXmJuicUmgVtwgxPq5g3mIQR
asJk/4SbZs/tzuY3ml206rdl4yxrVEWR/bOEtIOjRzgQOIw0rU3mSKdb9giNF1sRgQDofhzk1QDe
Q4W7wWxYLH8Tq4++QQ8aO/c4wH4Wf2DWroXQlomGQtJBNfNzRmB3fv8qEKy4wJvYCTBZzfRBkB8B
HXQ/TTOxtvR1QX5NMOikbecP7ZjHhqUPg7qXfuKaiYWvoQj5l44i8XPDckThUUJG1P+wEeNwT8Di
6GpqsGbUw8tx8r4JGYS06D4wcYEsoaN20PrS9Dd80NncTsjMvlZ+5+1DPwLjqz3+iAw4AVI0jMcT
jPPtrkRV24TqhSdBsiT2pr1pzbOTT08O5Gii4qGWXdD4W4hO+tEDkFGJs0DQBWSJRmnswVarCzP1
9XPd6t953dx6R6zF8s4m3AsauYymEAzhUU7jc/pp+jbwPE2LIw4i4ixrHzEsEgKKTOK8R25jO1UO
Hk1FVfZzEYYfrGInyQM+S48TgqikIQz5S4VW7sL1TkY5T25p4hQ7hsp8ezzyLdHrgdExqx7RtLUH
lNhQEOw4TrRi4iuE+iIp0PL9REsRJqlv0a34bQ3ORfRIJa/CoybMvngVAXzeY1Ghgryn103D7cyY
41oS9+0mQ57RAi/BGcD7gWdr3LtLrimJKFJmAEicGRSechPVP9Jx0XI6fkxkP+qjwMz+MzJmgFaQ
9WEm6yiY4rrkINHJk6JmpOPFWW2tLwNdZDjMy3vkRuTWLi6xMuWK4dbFzuwpPieLajWo7yCortk1
OqzB7mu+WsvDzyrU+MCkO1RW/AfZu13MNc8bJAiGg6HQwfBJvlo0X+tRXiDtJXAiAM/X7DiAwNw0
raBUgEtLKnEu9cm6+T4EAoP1jKkTRqwxIiQVVuYb7HMluqDZ0i2ujbZGBPjbPPfeO6fTeabnAYTd
T4eSLBhGAob1IpR26uq2U1lHXDqtwu9kP+1AM17Enym8YheNWlz2tHEAk2OaQwA9KCcU+7XxDOlF
AJiBTM/in05y0TSDIhhAOeH23hFc4aHYNQf4KWuoif8yIH/SSvVpJesK1iA6JJRysTE7KV7qrRYw
M9ZqyZIY7H8xhgbMTwC0zCpanzfW7ijURZkJqLyTBnlB4g3tLB3DpiMvXVLetJ2gwfAWhA4qVpOf
lF4+f/AZNOnWamx5NDg2ijUsoMSrnjETGDd3q1da2Pm+sNyKhuSZyuw2LPgDvSWKmyMQqLzzAhjW
+OlZvM1P+WQ6pkEHR6s6m1/lvzuzC2H7fDE5dqVwfHpZPbJbOpLQFi5NQpbFNifCnowxmnjCeQEZ
2OIqZ7plmC/MnTgETA3/7OazwfiFfJl7XV9bLx7uWnQfhBgMZFb4ghxRF5rdIuHU4ysWjPhbj7MF
iFKaRqPCmbU0kWZWl+fmQgvP7FAuDvwi8mKijhlWNvCdMV4hQn+Nr1PlG90h7Xi5QYl7rE3+KLg6
aJ6c4Pzqlg6qsUEl6cJvYJC/C2/1ghpTqe0Seisk5BjwM6B4wk97x0kZMT/QfOreZdmeTOmQaqGf
vGOPphG5b1TdW/FxrteP0FzdpzOkYhOJ0tqhK32lkBuSNkoLjUFRoFmh5Jlo6nt/ru6u4jY0Cpp5
cn0qn4nt1kn4nwMu0ZFRk8l6Fu1qV3f844uTmRR3HwhYesY19MEl13s3y7znXWvrTNpldymWJWgl
0Kedmu0aOHYfHDr0XbAGa5d8Bbfn4YIfT8NfIwr77c0dEHVlwe7xW9Ld5aPQaWXMtfRFw+i/Uxil
2BCu1otIVbs1pyu6xu0VZa2ROt6rLy81L7kA/zN0MbwxNp5sEYFNYQg7Mr/V9VUpLENYZxpi8+ZV
6XWeAhb66lK4RhfwujPMtLxd8sNesVnwv2Hx4XiveRhznJaeBLj3G5WsCzwaZTlXJV2+58Gyr1F6
f+qLOpWaBzHRW1lFADDJzRP3JRAtdRDaT7ymUSv1vDQrr97O4uXWY44pMbm8+g7y+umgGWgHE9pE
shiWmMg7LnTT32bLGFDGqrwjD9MZpOfiyLmDHoRCkZYbdQe0VboGsk/e9XXJBs2RVfxT7Uj2JIiM
hpZBfljctiS9zIs9j0iiYn+lDUv0DOQoRaQZhPZjEHR7m4Idl3/Fy3Yz9OdYpo4NvlavKxQCsGFz
2hn36cV42G7V/mzYHU7qaPtduNkd8dPTd50tjssBCOe9ut+hEGYyDpkj7ghh1n1sUSOQtCMyvb9t
WC6tS6/3MGzoEQ09SJfdNk344qERe/uf9Mp4onIi5KmHuA9zRpmVSNePpUHZIqfEgbI27bjd3H5P
H1PlyjSPo+7fTWtxiXyyGTNsDeKouuCYzLhXpd/dTTYoFI6PVs+gRqS2plU3BxpU1EFoBxdh05u+
xrA6i4Zv0zKZDzPn0qjNTf1+rPkI1dlQWwA6/9oiErteeG1kPu0yj6RxJBCWYHiSPodaJ/VTUwJi
2bLWdzj6FFhwf180Y8NTJvMukdAoIj/9jZv47zihSdyWUq0WcVY6n4EjS8BTCkzoSKA96ajcqcHn
yOX5oH7a1GnNGCt0uK4BjvHp5d6zjV16CNZ+jz4iuj3HvksOaIPg4qKHzeBGK8xlzNu6WFdc3738
9/YuoHp+3nfmZcRt5DNIavf7muDHtl9e4x4FWckCCYDPGDWf2X7NSqMM29ipHNtSouT9lMr0Cb5h
li9mTZk62u4IeAy5lKGCG2dqeCSVAbvbEnWLxfEGPZ3/hhVza6x4Wvyg1JlPl/gT8sDf8BsKlUvS
xQuWGo7f0M+c+kI1BZ+eu6IpBqeAAHiSfywgzkTkkId4zxpI/e5lPs9WZS1ZGJ2DnQKhDPfs+VNS
OsF7aCfhc2CQ4MjQ4yQqcjWuJv35EEM55n6ZQzVbsyX71eplkeTx+O8VbWrIe64+YFD0qyR+wt5W
HUzbIhkTUMpqt/THyBEXrfYpKwucXVStksJmRa1e6Ohqve/ZMaC3IGW1nI72/AeZZAR5z4RXuOAh
UCHn3g87ezCabk02OQDGtDK9xr1Gg799qC9S/L+HDbptfdTeHR2MCVgDv4GpnuXXU5ewdc4/8AuP
7fN+YsyKzF2iA8HFVaNIGuFr/CDzYH5pVnIX4vqqfEVzQOf6LyU+yfiSxoh9gIGJ0K2QzAEsnObN
i9+OQlOO4t6ZbVtXITo1RfQKDJbp867jmsu4XCRWYpclvZe2azYlLfU1uK6BkE3LyAGeQT67rLHS
csjzWwkdNsB4I3cBXvzmlTpbYT2zr62cLZDeLR/LU/4BmwVZRonw12w1VYngtwLBDPeooPyQ+J1i
PDouiq7Y3MmhiwKUmWDgOqA9se50SMRAENFfqLKA8axEZ1x3JmEUXi1POou2dQUou2EytaBZudEh
5l9iLxeITp0Vkvt2DanwZBX5LAv+sHoLezVQkYd+6vOZ3Nwene0h9wLEwzZ/KzrqtCFdjsj+VPlR
MwNz271GMd6ak295sKW0WYVcjlLsJHs6lS+vB76Zp5h1wExCx0F/S4FmSSIFGYS2EwLR+QdsfKFp
bdiFN4Xu7MZuSCtl8qcv4dTss3Y3X6qQU0t6QeBrqscT0rOXeatufdDie3B2sIQ0KA0Bh3ODJ5wO
Q7KNWd/a3c94W4ZDMTAMv4UZoXSdEnohVhj+/mZMwPUPfIUL/sBXoh7grNeMJsJiJpkQKMHHj193
Y0+qsUAKwVc1sIpddiiT03RcZRIJqx7QEqOjsuaqcyH/1v9lAwU4gUYdo+OMLd6R5yEVR5GwA58i
Fl63ighBGx/xSVHaR709e5EUur2X5v71/m451kChfgezL4L/VWaLs7f0uzvDhiqyioHfmhHNdXUw
gpkajEoWIxiFlqw6MXhCPCB7/hV/319qF82OPnqVUd86ZrNgm/zVgGbI43Dxem4SJ1MZuf5V58je
pT5SjenfAXfmdx+CtDPMz99Z3RrC68k0nT16TSwlnwElr0CWsBujAjoTZCTBb53NpAVBqz88dxJc
uHcn/uDPDTk+mYrmdZvPdm91NhZusj90TSonCQ9B5xv3DPU4/LoULp42ynaQlUh05gy9a+Ms3iRT
OSeeAtxYBXOo5mYsvidzBoqVOjMIsh+qWVwlQ96woFId/4VK0B8vUVYIVzJ4EEVl44kKH/zZuhlU
jacg0oHRQ1vBfsTmiPHy+QXSl6zNr1AkxdWeRkszEjZiJpz6lSq7G+CMEGnjmo3XdfnSRnZCGUdG
xeKJ4xGIC+FgBKCNDcuR55Nz5ltSNMR0IaAKAf2/dx/K9wcK85V/dZEg+ZWWgfr0ysDDTDuFS0C6
ZlUAjhzX5wrGPru4SPOELT+ozX5ZE/0ieSCylV8Na8dXKWb3cTuY8HGnBp6lwaMPYwAjpJzGvDaU
t8wiaaD77nyNwy1jZ1zsjMMzmKlzXIaN/XkL0OViKbiVU5t/2NE4Khd7iWVBOBiuvI4HuV4ioLrH
5Si6JV0eT6sfeCx1/cWY/hz/lG1TZPUx7kCslaIakTjhSfdKwkmYjkO8NCjT0nz0NFvTz/8WEZLk
f8feyDiLwU6JhCMbetRJ9iryviXMFuJaHV+6C+bQcnC3yiLhxnNo73V0xg6prhmK66dW3ktlgaTz
aVMRfwrzelKbalyWccgRj0nXJIXfxGckARegph3uSsVvDKfVQTzpO1pqM9NTLE4Sfoid0nWCRFOU
LiFXpI48mGVaIbH2m1r4MZ5C8wZSrozeBE02535Ac4PN2ZVQUAbeHm1mYNa3Tk55YOuN0Yx/B565
q5BO+0BnTCcdIhzS7srVg+9pF9Nt/tcKkhr/mRHiEMRL0hE7w3H17z1NYfcJaxRY4UZm7CAFPLkW
+hifRKixBXMu+ps0jbjo37RsM/eXHujG1Sus+FoKg6wPm1P57i/9bShYbdT3M0+yvipVvIF00SEe
jkCh5rR5VAvKvoFshkqpTyUiTIAkcKMTeOD0l64QanLbKZngmBIoUbVzpxO+z2C1ZYPVqDMedBtp
FDk2NnxYmpgbkjNl0V83kKosgdVSTxU8nlqdv96oHK0YfYnDswuSm53FZk9sV5AUJHDf3krzjidl
4bnNNevz6rMHEmzNVFzmXTgirHg32KsR7zSoWVT/Qw8Rp70f8q2FIj3uGDOi8CG6s5ip4MVB0Nu3
yNwTd+YctwZvo2cjp6qSXmeu1R/Rx4b+HhNv14PwHJk/GW54pav64Z9pL8RpR6tAHF/7nZeuPMHo
CoRLmjA7MbyFyxnVciDsbNrPGpxWWuKcmI5vN09zSFnpDmbcs3rJieg0A78EnMWeKVXdrbzPkUe6
Qz4pthURIsC4hn3rp8lNcvBgGOCXaFi6kRGIqRFKT03sW5WUSwEJsyGJWDh+eMYmd26w9yyn+NPX
vEBjSbYeimKaIHAw5JgbkRbJRyqXjYAK7+S1dCyuGZPsppGgn7y5xZUglVClwFQpobGiH1nkMQXE
ywffvGNkxQtzpxmEm+RzKl6MY90GpBhLQcF0KyRFmCddt6DzU0fXhDnsPZ6xfYsLauwfXucPGAlq
1pbvr20i8/dihzFBFrl2Vl+HayqvKZMedr/FSOm7DdDbw2ZdBodACvw910catWZ2kEcGXHzeipG/
B22hVXneeXBns422sxuD9iW1Se/CXB77e9/VmjQ1rwJQGgt8tKhPT1NEnc7JM+OHCdtIvSy0g5fv
X2p69XnMTGmZ0qo9JJaennXkHbsGTFi6IYjwcIQHkjNA2inQwnM2GXXSoSk6xUhjIQFGugHhhjA0
WtLurloWtKAYOUJDTZ6XO797KJ64EoDGVidHE/Lixd1dfecPJQ+k4Y2XZhREYbhKeUuRl1XTjCl3
awWc80UT0pqyan6jkTUjBrHsvWx5vg1WVa4jYjxtfj+M1OJw3SZ1C2k4Sb3OmBZCGKfMfzN9IoLx
UPB9LUt9EH/JWoJbe1PZt2zCYfRVOmIXigRQD9cpv1HAm6+tipSzgAIfI2JCojqNjW6lI215VdIH
l0NKvHuqteah8+pcEXphWcjuQazj46iPH9Rwav10z/6mf3LZuwO8y/CX2Tmyks/hZ3dWIgFn2xn/
ZKJotm6lQjS9tLwC0lemH2qyf2VPvgLmDVR0JuU7o0Ym800/TTpmAuBHmfdwJDiEz5kZ2lD59lCA
Ocr7IVJt0xTkCGKi7/ukXGLQNUOLYki8NTu4OR270v0cacoJF5ilfeLOVx0bK80/XpGfArm3h6bJ
arN6tX0QA7orNYeWuv0W8DpR/YSr/LTqdh1XAbr/MIbyTHfeRAmpT7AOV5wudNDmw7iiuWiFfm/Z
xqVuTHFdzEGxUlB7CUrLVRSZm+vIGzmIVn9ZiViNZb3TEdD4N8YjL7UOM4adC2Hs7yoWC7cQYXv5
swsBWSr6AWIxX2gzLxzeV/ippxW3mfUcmUlf/iX99B/H5I1lhgxbAbWAdoo4+FzUQGRSXN+KROgS
nlEYks5Oyoqjgx5nmF/zjkabMNBc5BxGxcAg/BAAYiphkGdLz2mcPe/x3gdlsas+8Ct0UyXkNqnG
JSb8vf2GjwHhnFFkBScJ8jYpBbK47hdZzgiHfWb/XXIBGJD+mzQxjJwUMkwaX24knES6cvWLKJnz
IcwK0+w3D6BYZgmSPmKKyBJNChjL9sTgWqWVelh9HuD43//Vt9Ym4KVFuT3vWCgR5ShJ6wvofKmn
TY3/kKvkQihw/rH9M+I/ggxwiw3caHUCeNbSk9LAVfjb0DelDcS2Oasqrvs79nJG+2I0kKVBILza
87vCtBFLfyhq/2OBWsGS0O3HnIY6PUROR+/sOUYd8x5T74WFU0A0OaDAOvGV7vn4QPc4fJZp/AyY
S419RZdRoIuEZt6kb1q9OpjaS6F70tEyY62+gdEUd11jr12VjQ52s5a2o7HRGSMTeCCnbl8OdRMp
Zi1Bn3XH1Y/WCuI2d6CG98AreL7NYaXUEBTmOnObsm2FdkDaGGkaDhzErlahl0vbivtdnGZJiwmr
eF8pj8rlMQNA9aOt3BDEKxNfbytJRwpdLHeVPYDCWX53BY5LyKSquu893r6TTUitowRRQeujxf+n
j9doA9dh1ZjDGAzhC1OO9Y/tvphS2aDFyBeIpjPEE0e2FFBT5DxAjGeFF75M0Rg8NqbCRxbCHPOA
FVhApfeenUTmsgmTKbLwWVZxvi/eXKu7pPc6+yy1kohsJn+kipLtsFZVoh9PLHaCQ04Bt+6kxr8W
uy6S8HavnlJD5ZmetOBTuJ9WX67WH51OacuBe50ghXJSRfayAfpSUYZwnPeFFcnQq81ppgYFJ8h9
mMeRJ/L/S6nBD8z/GJ1QwuF+VOky3sOprEzc9xB0MQsVJivMP+kj28UU/eTZSgUPOFf9ULrwmUeY
doBlyiPPSG6K6dMkkZDIPBQdlFXL7xuwoUiOMsY3ijqGtgxf+r5HYhvKGiCAwCKvlArFRbKcnIUX
UAd/S4bGvNnT3L3v2/+e3i/+SkMenOo1GpvruO0VfmMK2BVk2BgzwxAtOGuSKL2G07jIA0xaB8eJ
7P3XY0zaaE7BjeU2g8XU4dVQFjYhTMX/Fy0L7C55yyZsFOF3n+LFZZaKpPD+CQ0FfLHU8E2jBg8c
QW4qS3CH0X3gQma1vHCZSHph/NIcNlfsfUt+7zgTZQFK97Ko6TsX4d7xDjU/ehir5CGMF3BQ8UuV
RIcLlvAPam6EPXwuqSdTrXfs0u9rPdowar71Q45blvleLwDWz6dGvfc85qouXTvedbdMnOJUZd3x
0nWpHa6hRlRauJltu6ImraZDjiLNUR5I9xmH2a/1yWfCGx5qwRH284kNqoZMMpEbFEM6S13pCLgU
q5q02NjmeGHkT/4jWGqt6Ncyss3zDbbmdYVXMl1YsQAHOVTM4QXLQa5E2zgrC3GcmiB1PN+SjX03
VYnsER0W1GuIV0hr+j6hiPVwBHwOHCt/QSM4EpMcBe/Eo5heo+ZE83DLJvwQvLlyONr0MY92eVD+
m4iMVL6weY35eZdjze5dXUowzkTZIlSWNE9y86Xq2UH/NIkaAMGBT/Y0CLim0pmnFdRmuuxFndsj
vUyfaS/dTy1WDhz9mCp7daT52UIf/NpJ3xenhzLaaMQB4H2I5yYrfWCEwBhGgZKMaCWuH1lYYLXl
00MKJovJcOtGQo5XZeKpObs1jySq4i5SKPHloln85zzd56iaeugWg2gWVne1MHtfnvBGssnXP3o+
3/nEJuEQJyeVLk6cfVwsBBHWmK14v6suyYu2KVKhO04jjEno81AjhoYmP+ASqs5e2dPYuYvmcd5s
I95OeN+8oHfg1evIoL1CoGXjPDopR5aAn0T5wz3v8vDURgd5M2jI4+zJ7YBOS9XA864G5Y2hTvDp
h3SAO+qJ2zthWJQjclvhzVIgkM9ej7KUDreP+j/ivOiendZC9haErPBpIYXsNl5nnOdHE0mVXbM0
t8h3OtEmI4YgsND28KLy7JgtWhtZWcxg4Go7C/l4IMzxhtTzXsiOHCxxlV7rZvsSINcbKxJ3Hieh
rCegdr2KejETpUkCB7Nr5rG75H2M3gUAPyva55WvVvtyMfDbZ76lbbcgVTmIjGds5j5GK4j4g0Ce
L6dPUi6Mfywdh4FR6U0Xtow6OnMKWLTEC22APQL/C3PzrVo78v33shHn4qjZWiWInCZU8nBksgRX
RSOOn71fuj1KEMMoWxXDI+X52bj/EZSkMZgf0sugG9KQlHaVagWrPc/u2FFW/GXKzyk9u9C+Ss4D
94qJd5D3Km9YKU/lUrVfMbOq53mNw18OmKbIafML2PoSxdAZniHtApd5hTXrKfGC1AX14VcESykA
pgMfXAf0AmRXWTjpC5WWAsOfUxFQn7uEDt2PlinUeuoz1p7zKvwdRObFz1U1OuvbSzhW8NKZ83Wx
rFUl1Qbkj/b3x+nGWMU8npUZihXR0/KJcs4lAoBxuQ4tkXaszBlaYrGEsh6mBvpSaeNDCuw9QUw1
hnUpPsno2VmnzVQxKvOa/jrPwDeMTQIRJ5P9/XsFqTbxGRh9csOyn4pvr/v9g/VBe+RafjZbqr0b
pTdEgypT9aNvlhRHkoOlCheW8ht9GlUNeS8zDgdVDZghCwGnXXqWq+C+ecoSjYn5NReTPdZFwkxE
cKsRDsTqIIBJYXT3f6KqoMprkVCgNPW5I0LSJOATHys6o+z5liG/71fHVN/VLDGRaS887yFYgOFq
K/ftFNSzt6Q1zuxAP893kcZxlObK4XSiMxNW4q+ui9Qd1KMuDd8fMnLfe8QsZjjqqlJEmV6D4I9U
XA+NPbiqrDdBfZpUVZetEWKfeHjy1/8BoVOG9h0jpwb9KGThX6tbKHvVgK8fbmSPzL0AD68Riinq
uqv43nxBICZ7tk4cGZiSI6qARpno7czfI70v3gS3IJnV4nOXmDNQa1Fagpn3qGpdGpPk1T6X7yGf
ZuGQRGn+gLER1Y3NV9Y4Gh/y0rKWrG2HfbM29u3a8g050ftBvHWayD1KlIC9bAEw5mrBWVy+rRNk
MWyl/+J5tzKNg8OKD8RhvQLVQrSEiWPYepcR/SZPDEszhYAIlIM4r3glQnf7XRdOf8E0fewciV/G
Ozt0qwYOLr21wnGZwsPgWa2i0UlUXOwuz+LXwCnPelHkC9/ZrpTgsDZW/SlHrHmNxWRAx314j6ne
tam7cyE61piH6UdCTQa88tdA6iQtEnAo6fOFEplM/9+nSN0tChT86BpLI+16ub2LkvtNfI5rX2nz
8TW9GfVyOxipGxUzWQBqn9U249mS6fH4MFFkyifvgVyqWYhCKL04CkPZPHQh09Wp8EyC8NAyTC+n
ifUoQ/cQCWyuKNbHIA0wSo54c1ec4Hrb7V/F+ZItdwWjE5K2wXk6JjGCsfl5BFta1QsTT0W9Neck
MZCLsV2xhqKtqIOX/1em7hafDBl0rW/gpKqs9k3szmitrDLOOCzqFpcl6M5KrqrJKGbh/+hHtkE9
5XdzVTw1LeK9k7ck/6gcuhyWHkA8K917jlKxj6lTxp9cf/tEL57fz8gWdbcD+Qcgzm32g48aCJr7
dNUS18lXrNu1rRVvfVZbrAR+hkYTABvC/Fc8ayGgyuAD94pQdU2nbFkzbuXDfiL74ZcXGD9pWCfT
vzk+rp3+yEcYw9vDskeVrIsM0G7TpHd7bdafcLLK6Cmht4qLCShpMUeAzlWZJngmlopqNEBqZcDo
PajrzgrLsJN0KMzyPaFCP7BFArWbBnOGNW85xGtiExkexQN88z74So3JKbtB9XDzDT607mNQKBya
WaK0qXA2TdA+MFHAEbUAJvHNTtIflL1rfjgbZiZNK/b1OyPTK/8BsrOVp9OSEtAuagTorv+D791j
G+4RPKs2tCaKeTodgLOt1i4fpNvBuHCLm5IrTi+bAycMxj6Rs+uID8QF/YfUR+S5fSeuBsDtNNyT
kyfQITz4J8pyfgh2oLDPTysa3abrlIt8eIPNm51CuqVzf18FJ0Sb8NYneWGfCIZKUZ15oTG7tImg
ZPedY4pW9YiECLUooQ8HBsck6o7NTT5DhewIf7aoRIL3MVuBAFtKNs2miBTRS3+7cFkmhWCD3UZo
SUbRY9qVX2AsSdGS5Lf7GeRPLE7UUqt6FW23P/z5P6CEI0hgvUXkH8JvpmNVTAuGrFAFivYA9FSq
RUej+b21Erm3iZwBb+DpARms4o0FSJuNMxRPJa4286nro5TrAYpkQNYTz8CjbplbTTI9h4uP4eAB
5Fmcl/PTHVp5zVtRZ9/7US21yNsEDCWs1U4DUiZBc7LoOa0fDS0SolsbS/ahj4PAerGwoIZe9q1Z
FNmbO1niSlO9U8TUEm/SIvEV16PJCP5KuDdftoR6CEGk0dUJG6A/bjVok68FhwXo/MhwBSp0itGC
l/4l1V6SG2SlhBoJIMVeFNO8WoK14MQgUpNQZVRNxC6ZwWvrfCrbaa7cYwTwDeoWcpUoGXOPVCJA
bqcKl3wxiESgd/aJ+E9IEhSxkEdB8LJJZrJ/Ucmla96RZxoNalfLYdIY48ZNw9f+fwlaS8+arat5
zhceVjSXErZb1quEZMrc1sS1wVdfa4PMsa9gAzDjWbGplcenAoEc+rMd1HfhyLwi4UeRQu36e1a2
cBAXiwnEXrZ4fU4RI/MZ1mBTkSeu9draraVcLoLvUg3xa7API65jzKdyrRXn/Wpjhv6JeI/WSZXB
AVHL7H4eWLkmu5kDv9spVMYSw5rbU0ELGJcmKpcCNa4Cp43xGiC51bN+uo33RZn+meM9ShpSAbsg
cswJUU1iMR213ohTc6cehzeE9xKCwi4+nTPIMbS+/QyIOD7OYLFe4Mlg+drSG3O0bB65CRLe48sI
MmUSPU7Dd0n7oSrQyJVVUymsCOT+Swvu+NwrgMsXCch/gBhoZGJ0kYR3Zt1JdHl+LTETMTsoRzJd
IbnDn0jeHRMhP8sYXsJ+qYWQf79doeZtAkpp6PKHMBXPw5BedzTFTlNMiERbJ1HCLfOANs9Z2h8C
uNzkbd+qvMxT85pKZ6Y1rdA+XJkHI2tJRZw2O8bw+jidB2330h2P0lYQWWOpfFn/Kz9YguMZGrf1
gIGbTI3Wlt1+i5uFc28M4RWSvmbq3ouRnc8XmfM83apP22XmzR7OIcfXWSUbcBt2Qdyc2Y6ZI7Sc
1eCj4+9vGfGIQUfMAnkCmhCldl9ZlKExrzakD7RpdCRKY91FyzLtjzoi7Zsqh2X21+kI4ubaRVT5
blt6ma5MIDUoauw9pz7nHyZckOyncwH9xzOgpR6hqVPKa0x2UbYIgp8fjQGORblS5lVT9EtQFcFZ
lfc6RzGzb3WuUm0dTCsaHlezs62OFzugLRIomnnX2ITtoevMUHJsgEkMADCo/geRwXK/7cdETTVd
X3y/DeHaYpYR++ykkT81RSCtqtFIxbPp6nvrr/zxm3xsuwWrQ8usX7vaRIjlSdLR0LwEzSdDMaBf
Z0rV6TdSepm1Ij2ryNY6EEMyNxXoDiD82fffrJKqmnXPaX1XmD4e4YK2OySk1SsUo1cTMlUjMwr0
j9IoqkYhIzuGtgz/dIiLf0A64GSBn39jcdRiGo5wxMwcM4q4PvrhhcE4uilpVbaSLz2Im5arx/6k
7cB3Gkiu5w1Fp2yts8Q2O5h+JBP7c+jm7BMc0lim7UGBnXQegmNwGevBNNH6nH71AaAlNel2MLru
Jk/VLXkSWakN56CyYoJcwU3loRX2thfrcnCDPOzzLFYwZotA2rG4O9IeGxQy1oeqf2VuormH3/FY
IQCnSQkRpVWJplolDGNKtkCG06TfXVMSjeIH63Srk8LVvCMkk5RLlaM7TN2Hi6mSlvnvkP5NBwBo
Yo1J5lNgI3npHISEJ1/JIJilx697dOYz+9EtEfoxqHhGMSvsbVM3IBa5uUibrgJDnnP3I7FAqsAp
/HQh6ThlV7/faOPgbzv/3INJf0u6LlS8TYxT28qiCDoLsi6De87x/MOvP3nXV6q5CEl1YpsH1VCS
t7eq+pOf2ItaQYfCaNQh+wV0MGjbQzlncmaUiPAr3ZwW2CUvdwqg21ltsNEfLK+MEcmeo5KGRxqX
Em8AwFz5uf/Sh1MSSzhl1ymLAMPxD+Eiz1uTVJm7q9edpBklzlQ3HyJkA8ESNkqaV+b7FJoSAZxb
UrvK4PgjN/UDFI6JVxNrXHvhZDqrAqRGPf5ejHTA+lR/qYl0JahNHg4iiet6MYsJafLXfo96vYWr
e1nVA/Y6yQM4MdWu7Mmyz1GpjOtdKcYzqyK/UoIAQ23470mszkQIdCQ+5/jq4UrU3GrBLbTqW0U9
MAQ8LHEwRopzXtVFH4o4Eug/8VkkA3pDUUeDhIAPz+9kAbFGdfV4gO8yELOkqN9YdFnyxbifX+na
Wu/weFd9YJu5qimKxQ+6O2cKQX+qgadJ4uAqNj27DSLWhizvnqkxCr6gZ/pym+GB7kY2qVx8PyTt
l6cb+XggZc4htAY1DsUSZRhCfJBL/3NIw67av12DuHp3dXnIt9gDRnq3XjMmb2aw88EFTFbDxy38
W6OHM/rOotWs88mO/FCtXgR+W3rMYk56jAeTVL1/bqYsfPHsBpIHUvwI5CzK5taXSzZBUWtbdTDp
n4pXAS4oL1NF/53FylhAUpSQxXPq4acwRMmX6LkvwbWDKz0ZcrkQDBSsn4p+ApxwI6QDKleaxymh
jEC+9bj7/OKGbg0fRE/puWuoxA/uTeP5A/+gu9VHI09IhGsu8TQwAXecLSMu41MHpV4Qev70zOq6
x5Zzqa34/LXxOOuzSNST2ikpOIdKvwnqYHTn5v4gXAFDEgCCqR8ZYMrrHp+xB85Lsev/Z/9MqVXp
C3qgtuDL6lY2l0MLZbX2xlTdz75jtN8pxUKINVXEPNf7HGphrRxJhiYul9akpzhlPc+rGsPoEtdx
PbFtPxHQQug1TEbDSadlLJ6lBFvNxYeYwKi9lknfXu3UsdwBZVs7GANc1F+zon6womS3YkalEhCB
OfBkRrdTOmgJkVXQvxi7MGoJ2tlkvxBKirAz5Me77Wy7XcZJ8IoVZBjb09/wfvCRdxDvGY9T7dVJ
g3+bUTeAaEMdyyoWCR/xv3nsFB2djky6/GlpxdacIKsVTMTS+eGljSMAZxcyM9ZdgLhLRWRSnG2K
eOj6rPhD88TaC0AT6/c2X7TO0r14jQRmeKrgv5u79j2azc5zEFCvKuaYr2bCah0N0Y9gPLSfMqRM
rp61p8ew8AbWP9OAlDKMmRLR45mhASStPnCCYI0FkzPS3MTys+jiYxsuCBQdddO+7BnSQFenw8BS
jl9P9br1+ZpQb2kElmqK55nDRUu7Q6MH0M8vV/Mm2YquVVm8oLZ6MlurfypQexyqdfmLiL7wup+g
JQ+djdmRH2LhDV65vbSzY/amSxrQv7gHOWV16PGtg8Eo+nU78KndivBhS18APiK8QhVCundCnTUI
mOFBPwtDbwYenM7754lLrBl8+bRnooltFxA0N2H+bnlntoI+tSI+Eh+aW5ZXruzYJKaE0duHAPlC
SaYBVLDOZNkieriA1oSN5Fk4bUOJGLaNWXlk/dEn+ZVMwLdJN7xedWncGesixWSTpnguEG12UGtW
vBuhLZFwrMW8p7kRm/H9bF4fdW/jNzMlarK1yzMw4qJZRUeesnadRE0RP/K437zFB5gcUIvNSkQK
HNIYlH2G+Q1xTT208quX0MZ0tdAJGFT3qPTDi/HNvx3696gXvBq+PCXq7yLKk5eeSKBV8swfjftR
bGQWzPZNiSVKJBal39ihdjPsrHCioSaooDdcL3byqNkVg1yjo0hq1ws8oBIt36HkCR4qnDqtt9Y8
j68cGUHI60Y/4AHiOgnXUBnITF8/CySABbIx0Cn5YjBLCl8JF/w4YBsbDwycFNP2TIrbTGnU2mx4
cpep4FlKtPBFgIp8BUYICG0fF+E6eFnrjNA2xHZnwLhSFtgtEYDM1OgADQsgFxRxKpDbinVKnLLU
UKcpx5Ny73E9ZqZP9lRz+2xtADnRaiUXbj3q0IwEj4XhKdEz7CNaFQE0bkxErpVFRbeyrJJsytxc
BWqdjYzRcT5SPcASJBfc9w9KWlgI4rdrCTtUa6CCEKlRPEIAISV8dxyUOvX50c3YzaFnLWaPyaQG
Zrv+fWEaWajzhSH3XFF8/ZTvgZSO9k9YBQAx5XyDjhE8R2/KgwaBw2j36VWlPTLRukoRs56bQ2L7
/KhsSajP6w7XAaSJZzLFDWFN4p6XicMyE/pNLJ/8w9ZpfeyE3wxJm0ciwq+T9ZT32yrM86bP9mo1
hGuphcE6eyjxhY6RB0tM1nMWQ4y0A6pubCHfl78NF1ZO0jTY6WQKFgCQo4w3ukKoOifc96Xvz/2s
i+vOUOJnhqVM3jH9O2lbvJqwmTO4wnej3PFi48tw5qpNLoXfNmxjoAmA6VxPWS8dEK9qOtolp0yN
pukLvn1hX3S9Cfa1r2YXEl9l8fErm5c7asLRaWwkgrAi8QHr5vqim7OLQONtFlq6wAnfu7pqqKZJ
Q7YYIQGEmC5pslllpB7RZKEUyxZrSnL8UXalV12vs/9nocHn6dbWy+8IpH0Sb0O3z6jrbPdQbIWF
XrbRUjU5WJefkV2e3mfj4UsvyzI1Wqsgvvw0OFLe5DgbfsOjQUipmDRod4+bLXbmsS0ZgmAq4eH7
Pt4LZSw2PwU6En2V9yqCJqFcs+t+xStI/1o1wJ4oM6j2Vl2oTBprzUPsP5qbtUuI+3reLBNa8UFS
vrtrSPSwilXYJnKED5Jg65ywhMKKsKvB3ymzGfzPhGbD6Zqu+S2jp05zXKUOSI6RJHrYqnWHNILJ
hICzNYxWn3lnaBEKvATBUMUSqt/uIsphzB4GOXr7Dm348mMtQ2mtM5adYCP/C9NKyCSFpKJmpaEI
5T+vTyvYeAuFNQdgeF+3ahvCKsTcdY3zJvnh9Cn5HCdYIqMFZ8c0Bzlw2nOANXCzb84FQy7C/ft/
4bPpOy3YI8BRUTJbSUx7ka94dyHK4F0n0FSy79IAiw/t7DL71BSMJ9jkgxry6tD7j6F2/L/Sswz3
+PiSOatiUFyBjjepsqUmQWPqdBl1TWgcqUzQ7XMBWQgv2PTAthKXxYXXky6f11YhQs1k0whhBccK
q3wz1iXNp+qsfugpxyMsB8bYOIUhD5Dur1/1xAmsMk9PE21UOkbGxUrkQnntNOcrTjEUZK3gYsr6
vTZ6mIyTMPK01I47JnJQx9EoioTK4zkErfHRoC/Uovh+ut9k3Xj/mG/WO8i/HJwAeXUgn46Ul99o
vT57ok0MxtyKGkVknHPbx68LtHY/cvQM4RePpo9y+ceNC60DyKoN+6bRknccQCSYUZ+pDLH4mE7P
/P/VK9mMH63bXNAVgntUNSTffJaM7IEOnN6gpD6oWGOd7MHYDgBNUgLWByB7Foqt+h1uwTlC7I1A
Jwdpm5JEdWY3mYBPdAh/clX6mh6tgg5OJkUlVf+LrfP4P2vvV7LQpP+4TO9CdgLZMRHBIoUcUQzK
EJJvCJtJmsrRePMbfgXAXHh77Puqr50lki1j1wr7Qa9MNCdnE0wVwu5kPylu7jpdurGq8gKN+4JH
eIbLkMfRkE9Agf6mp+h2ESvwDPwWoo3iMK83U7R9kLCphXUXPqk4i0beDfWz+Kmck5h3S+5uZspG
jL0QRQ6e/2aFECsvgHQ4DIA/RVQg3yvLgzMTN2B0ye7VP5/3os0GsZRvet4PiEuJTl+OUNGXTlQG
u1LSc+vGlmNMlcRwTj0j3xxFGLjY/f8hJitIGSNeUyosPOguWfifrPF67EEvxBnaIo0IH3FG40J5
fgKY7FuFx/LnvYvQkbPXIv1PGfIYdSIqY/5+b5oo8LA1LXfyF6PA/4uBlk0r98tBqQLfZbaWSAmF
bm40obnQ20yFo58KnPKiqLSUzDs4qu3AFMsEfT748HFdolfUzZDcO7JRlgtY9rstVZg+t2obSWAF
TuqCcKdT9EzNn8YldJ6q6ZXogbEBcCYQjYJnjhRPegwenvBN4+d/qCfscjO5WfiAATtej3m2pWMf
HvmMKxsJW77NWrVRR+l7mvpqjT5aa24Nrp6saSLAf2FdhruW9iiIY+qlV8Eh4H859d4BufLr39wr
XJyItm5I10dWuVmS7XLvlyAzog0H1ekEDieXJCeblIPj8NynUzWAHF3qT0+KhVcBybZEJJRNyQEC
FJinlp1yikI0PQQZihK277/YRbjRYDI2kPMfPl5cZOoLf051kx/iBWI4MV8/P/xC+WvbUz/yCfLM
07RqLBppXfvIBHcvdjDzn9fUIZEMHgwIy1L5ac2fd8PdQjmh3bap9/oGpW5prTQHQcA0+wKz8752
w8wkJ/NpQ4ld8PN1PKSqjt8l/lWD+TFSZrwye4q+w6QY8MPZ1AiTGA10oKO5trlEIFUlnlZqDg8g
TXSrrl40230236xoH2UiQSzlcLKZp6MdAXPQWx6TJcQ2irGkXHETb7+feEoLNRI3dNCduEH0X5w+
/GDvpmfxyJ/o3KV2QnLGgiP37r37dPpWFgjDzClYWaZRIFLdXNitGhcWXG/iVCtL99XPrS5MqDdi
NAqgRewD0/KgrY9r6qWHks3UcbQg7d9LfPziboEu7+/X2rL1fyETi+XzPiTiZ9ENEFEcTlks5/dc
xxfLoL31oWVybGeyI+PFB5V7LO4Q9Ulodof93zkzStpSU6ruxdEWnb6zRjQkh4dZD3eqzaI9qc2j
penRFueZ/sFDTB/saW5Nv2BzTWUGQChAvpdJ+l+eK1VDcbc88FTTCXMYRJRzRuMtF/QBBagFTrSm
n+pg/GuiBmeCDaCFjcfCQ+jyl+BOK3YEgwjR5N3DHJwMDgG6Lae/W5C2gNJp6Z1u80B/tZb3WXzW
uHhwf1uJ4muBP1KWWlYTxJw8krLXQvj8sVmCAplhDwTTn5Uq4U7xbgRETUZgCGhXsdkmmscU4DhH
0Bw3mfP8BZZdgaMtJ5Km+MrMuYK7poZiqpG5XgW0KEMXCwqxZGnD8ppknn8FXgzqH9REdexUzlDk
l0TGk4TZW1BvB6zC7WTqzsh1MePkNFu4U3QE7j1bvPQK0acaGuUOSCdaS8Ow9dMVqyJhwGu2ft83
A3oS5nMxu4+Di3s9ibGquQe52UKSi6t6UlQ9yGj7rUb8/XzXWzBoDLAufcwwwINWzTRY0zuXVFeg
Mmy1gIc2S3ytumYvo53iRnVmqTzl4OYG6HI8OrfkqscXMKsULlCm+XBIP8Pj8awGxCOhBOfr4VCT
kHDb6ZvNROMZ2574rU1v6ZzQlZc14s2pbkeKehNzfCjcxp+JeiRPoW4GP4oOJdu/pkKRagSsLkBh
geIchueWboQnnjfcomr/5usPNjNfEnEDKnTQJN1rwfb0WFv4ObhDVaiRzTXMLAgnbUD5mGciMOLR
4vCxcSbbVT/WhYmO01pf3wSNXj1Gl1w2qovPko8tKts/CpkD1VAXcn7sRwpx2JK7tpaxvjvajmvF
OSia1RI10frJnrrfvTgZ5jeAXDESDGRE6xv00z2lxfnpADcU0kvwdCCpmhVbIoSt86elMp8/RzqD
QcPTQvc5VSC4TVM2Zz+AytJAbm4BLFI+FJFTmNfXsf49KJWxNRmIaV5V6z6v/FaBaIR9twjjxI4r
O4VS3YtKTUPE1rDT4W2Ma1+zucUD/NcvYfV9Mo06pXLKBEJziPXemAM5Makn7tmiycV19ro4oWw/
AC417MVWTbo4PllHvXrOpL7wXXn/7TikgP4V2aw+Rzf+BkKkz7HQsPSIKwZURqLanekU8kT3Gjoj
lFunilzrDeOfwf170X4Y4eQshHVMt8wXKqg+YQ+sGtsfZWOKErdDxLYomaTsq24bAYVQRcKpF/S5
tvlttHojI3ZcmVRm+H+yRiMoz8ewyI1KoxhiOUQEIlArEejDZ/BUDy0hGJZQFf588nIZFJVku0Nu
IUFmaY7f/GedAiUk7SAg2MGxF8Ixys1EOBTMhGrN9sTuwNb0oksfB6ZeI4Bu6a2Jf2XJHE9Xe3hA
uARQS6TFfw++dNjM1gNcDL34WL46dimnsSA6W8zRDclIbzvSmsQ3rPiPlZx+nQgc7w++Ly9QSMU0
wuLCEnfj7tmMmhg0IOC8863pCqNHvHgkWCy/2kJ58R/8gSNalOCII2dvB1x9oyKW6YH3+gTwtQZH
Mo4UuYTQKxndcDRbmPXQIQU19aXggLuWThMDSjPcBQUO4HKPDKTpI2Cws1r9rPd8ReivrvB7zPgn
4B97PATVtST9B4c7Sci+FZYeY0FKoAAuKPj+NWB56iiEg8ELcC2m4/XIB9NdzJObWJxhC0STgrMA
XENjjDv0rRDzsfnJzcX1qhbSUWPdGFZk+k2t0cY9qY47zPXLRxylms5o7CDnoS/kZ+n11b+t30Xa
UnpX3m3F2A+ElMrBJmpYmS56JQROyU7/qPs3UUjXyKUQf26aDwz85tII7ahSHcjfuPZJWe8Dki/D
UiJkLMcX6HB5GVqHwTJ2dDw9vZwg3L4+PpUvQkXRcjEgODAgc5vQF5nOwgW9yUcGHDBPn1J7WcET
J5094fwovPSOZ5WitGV900MVP+nSE7aLWU6li6nuDPZ1rpmlFS2qWF9XC2DLsyok7nNcX9rDDMTG
8NLMa3lC+B6FcHDRKM43pVC3zzeO5Pvj+dmmD1f723lnPAjwywZK7T2l/bd3pUmAqWMmOVQyrbWm
rtbj6mDPsULRYqtT26ONF3Xr3SSmRGer4PkgKR0rbqTucMOf8E3Cjd/er1WPAsPP1OD+/gykW31/
EpRhoV4Xym2dz67I7YY2+YCzK/u4ULWaJFTPTSD3Ds6enao6YpyR5VVO3a/NKvmqmoimiVS3rJPv
KJdB+sM8uWepOQ7yD6VJOG670bdiEPShRJ3qI1KKoxMk5Nb9LMZsVEvNoOxH+JAeaHCDUUdl/9zp
7QdD2Xus+kl9SAjdx1Kj5cY4/i6OlTnDFq4D/Rr+2AlrQZvXZxP9ndS3LnMcpEYAExomtP2rItJo
MPgieMt7fHFhiSAuQhPGL+CjvKejg/BrDge5+Y64EYpgmur6JCIAlOjfx0wH2KnP43GT56VS/3OT
NCW+lsecC//pwzLyNlQu0dbq5bIlailKDe/Qs7X4DhR9l0bcI1qYm5mMVt8xY2qkM9BJcweSddnV
gBZlXm31qa4HKvlXw4hYUFh8XOjiqnf9yCZWyN6Y/FXItPMHDjV95ukE4S1NG28m2V4RxczpO+uG
N2ihctjsWKn6tXRTv8AIjpYOEPgK3EqAAML/RBoaqYlnR3Hh7yOWh2EJAXqaj6Hc61GA5D/vRsd6
Q/sTfl8XXKMH3tNGoyLqLgdmijyI3viaot35WAH7cv59AXEYTOI8C9KoVe6dwM1rOVuQjaHpUUTA
TGQByNQZt6BwUMNJXonRbsFK2Vt/qfVFjzboiylDQD9BbJgUGHh1QG4DFKtsZchACWin+RIiKlhN
1xpz0XeSaVt0+eXghXISErixvMbrjoPHx7Rs8+g5prq9kHgiZrufy3Kwnob9AjM6EGiAC5axPeYG
z8KDhemwHWcr3/MSsf/cL/NOMrVS7tSvPzLm5ddoaB4lbTghsYfEo9gp9Zc9J7v+dPKHtkZZIfRV
VI4PDoQdtiNyoEaS5FNKYZ15wOXAiY5HzIpfWAK3JktlCysddylYpzu2yie/olw16ue/TkhxSgAY
PPHR2NhU0lr7EtyTRXynxD0OisrTRcHWCdgnxxcmjbIqsuofKPn4ya08YcrBKvjYvWCqgubfXOJl
/wtBqcJ9EKKuVd8iZHBiciWcFOkYZGjorZHH+iClKNRvQC+ySMrBGFlplQmdsYXh8cR3hKt2Ud/I
uxO38oo37DhVd/o38WKbRRCsx2YaIa9EePJiJHlLgGIK8RppQPxsOuX8xm4q/azx5DtKgnPkNKfq
vo7GfhGfGzpTOFLwQX6feg5Dx6rGO4l155kkUrYGZINqJ0/7w7ZcyO8grrXgjr/lHKVwMNLOnx7V
JZjweDpnZqbAdjoEqrSa0Q+wpb8KHPygcbSFnVf7f0gXVMITeR7YvU/bSkbaMi3HDhpLuqDd2+cY
RcVkajMN9QwLpxHRKlsF0UT9QoVMd2n/32VRRdaEpUFDFOjACIT9N5VTHI/AXL9Nf/fXM0GOC0mk
+SwyaSiVzAungwtROZ3RCvo9htiy6xB8CF/e1SMHG5uSXiMx5ZMvqJgZUHBrFr2uj4NCvdmgZmDp
E2HjmMZ8hZWD1uJP+cvzNj1b1c/Xe1PQ/Epcr6kB2gVldl9UBTyj85YU61pBV9HbBlXE9igq7fVa
qomDNP7B7qRtjRp4PZKO9Gw1deVQSKCt3fnR0oCrN2WW0vP7pJEIr/x6i6CUZ7h7GRi0YRiZ6Fas
mMDtto4vWQAdPI1nz2cv55H37Mql25MTpnVejCtFHnF61bZi4iUUy7cfcJZaA7QShw4YdvefpBjd
ETVE11DlwUBz+7k/iCC9GQTa3NqHj2aXa+6GQ2BQLVkEYKPTR/6eeYjD2Lp5+a8RsNrLrXdVm7AC
3E8GhKJRlG7LrhYAxC6mxcJwMZPiqKzsKUwlCOiC5GwXZpaYfQQdhzMEXVfkd9AYBMlGXQ7R/K9V
r0r9N8fKYTzBJC09sEhylZS19//57WF8MxiydUe9IY+Y/kkSStA7YXqFIRse5/IGEyJ9G6ield5t
hvSb0sNPeq59W/C5rjVmkRQPHWwM4f3eJLeU3f9Rgem8VLhfVhsPftvPOdNvb8SP7qzAiQNUe+Oa
jyL3ZCw5luF7JjkxDN6Y03It4zq6UdhvI6hyniIfoZIOFVjg10MzZnlI+2r1hPyHaOjKXBrcnh/L
/xEC5rdDLBJV60pCyMrtV8yz2BP9lwzHUObXNtdgBHcSDRH8sMsqJVrVxdexW6EDMKd8/LmNxexE
u+3G+yu11ipZGhKrxuizqpQysHGPaKEeSHgWq45aJ+CMX7rtfbNc4szx0plHGt9aep2OX6miPyX0
efwYuCy8vEntVFpwk/eunqROjc01QF/4JPFCuczCGdRX7rEAiJCckpt1PdiaklQ18iqpMSY34Ikj
gebW0xhTyQb39riv74ggbJmmWfNnVG4t3S0CDM2SA5Gn7UpaPTOj6mG8ua/ZECUZwPwyH5W0a7Jq
TrERZVLkmbKEzBQ+kJzd6WwxpOJfbpeBti5MX3gqK1xckbrE5Kz+gEukIAccbj4PP9ywTq658xlr
1MYY3wtkjca3ekhDnhqcR54Vr+ihwCMUBOZ4Td2IIodBPFnm7iMcgkVdq+xsmDyuocuPCpukaasO
U0uQR3aCbNtitnYdC3riv55QGflLm+WZdZX3kU6N3c9w2wIO7amFekpDIC5QqFVV4SqtStnN1BsY
2W3F5x1/ck1AHm6zx4UdC0TtRehTXCgm85yghitv48nQ1gRwQkkvbJthuPxU7M6uw8qgP0b9UjMv
rXit9GlNTjmfrNmrdmAxHzykA/SfXOAkamev9yid+HPnoHzKdc7wHZ+ta4oT473mFHlK/GYv/8OE
O5fFu5uRlg9hWyEWXN9u3FC69crLXOX63F2Dhi9n5dP151q78HA75GYBVAQNcr/hFrO+IKUKR/JA
c1ljlbpgp2BNczDThDL535wb7oSD48ZIATLDehc0ARjHsT4jnU0Aum6Yw6vwbLC0k1KcloVng29L
3mygMUSS/kPOWF5JK9WNhwnJwAOPHTacWairUc7C8nC3oZv+6Nu6lGKlEwMoq+D/ew3XOnLzaHPG
o8cc4+qA0av2pmEHvQ4JLd2eQQwofAazmvNkjU5QPvfok1vsZEf1ndluuDc5ICwXeqUXy7r2rY7s
eJCyF4L/nfKzPmYFIP79XuE1hcO2eHAmWpnMNgvapA4JMfFcERqlPDlxZuW4mIORLh/W7S0c9pcX
1/h8Srtia3VPZS/eXDktGxFVZhUuVKTSjQNOPH7+v4ai3sQcs7+LBX5F9bTgdLSRhDiuajolBBfc
jhf0ZoDPvIgNGFl7eTUGG8NDK+jLjYPGv4BGjkn800eeiglRniiOqmne7SkmMKiUTKpZY9vPXllQ
8iufOpEUs7sRqdg+eKIlZMSGKyc3cUb65pqwaxeQF7N/tSlxnmoC/1YKOJAzXkC6cUL0Lkk8tNT6
8XXFvqiORXf43Slq9qLRGdzwgSSBSbKWvKsuzK7c17k/8WFXq30F4M04BjCQMYrs7JpjShju+fHy
Edlxqfvq9/Cim1L8qpq7OiHWsdsyo9RBjVQCtGA4PK/Rbtm7yPGe8HuQFbsD4Vo+gHDy6AwyzEiU
aAo2bKVu+hyyCW6j+WFnkUPXhlcTosA/Rfkgji6fYkIVOuIo5EQH3UUCuc1bcJIwJTzWHV4kVZfi
F1KhZWnJzHElCrU4qfsb/iJ6FCf/3D8jzTpO3ZHAbT/SUgXGn+zJLLAJBe3yF7yoKSQwXUnq3zDu
00sv0OQj49eZonQ54ED1UzLzyfNd+ANw9qk6/CiBO/17f/Tp7s9I4o1WlBX+IeLSCD6S4FW1NOnm
+SbjxReCbETQ2BAQYF0mcfSYNuZyOxBsMMQ8Fqbfc1qzHJsPm2Lxig/XrSkFFYgeQE9YBYJNkXae
VdUGID52LacTRbX+4NxRMZ/Cwy2Er4cjoPH60nPUb7rX3D625MuwufoIGjoT0x/OuVFA0u8+fGr+
TjsKz9dHsY1qFtHGu/gL1lJoLJir283l1TJenob4GoA2MdxKg+J8xYGcv7FM2Gho7M1GmhKDbQTx
s235Dk+hvoDbn0b2cgaXtLdM+v5W8TRY3rqWg5nLTDfiX6EuX2W2li2i//e/WvpaVerADx4C990q
6Jbbw44E2PoTWZX0LUBpyO3tKRRDURqJdbpSaBl2wy6xGLHJGxfYm3TFv18N1qRb43AXjYQPT9aR
RZOa/uq6v0xVgNWTyRb47CQwRSF/dT2OeyCqvSbR7J4pKd/KZolzvuhR7xz5iOQ3rsrmhM3tQxN+
/Y13ZIBRW/dSf/G2TV1kVz/N9UhaC7CCmgZVmUBeJcK1wfVF2TA20D/C69vvJgdvraI1Y8k1ZLtW
1BwtTuR8SfGNHYaCHEYjcqmGcguC51wFSeP+8CwzE1ueiydj7e9XnmeY7lr2QOIGXmwlYd2AGS58
CVh7xp8d7vXEyflNPdIPxSlZgI9ju1gVXR13VyzTmZMO0hFu7YlyHtWSkzhclPQzAYp/yu5b5D33
zqSB3YnAxG2uzDKHTq1UfTT+3lMKTe6R6hvTfZYlo/pos9EXaRuRv50RiWn05vqgw9WUr7TPhHX4
oa8bQgvmrCwEtQvL2K4VkuU678yO3vAeVtCEVT0qOjUPSBioNmyCt+iyAcUQbJZoMob9+XWnl8YL
7ya1HiWt32CaktRFLNWgeBpLwrUNS+nxNir9HFRW0yuF8faUo0bem8Ws9rK5nETydKGNyY2uzri3
iHviNO1hjHDZmpyIHn/4tVw7xao9ubE2lo14Z8mBd6yp7m1KctoiGIZvHs4ql6A+//eGSIQcy7wx
1n5KkBulixqLs/sw+FB+OYxRCn43IYr0YwNo0ig98TZ1AV+l5a9dGOPEFHKMnWuwEfJsjQDCsoLz
6IIldE7MjWdKBB+VZ5S0AOu2cAD8mZx2ZPfTefltngqYNDKGKa96aEPqcNfORare8+YDlo9sRJ+H
YSENxOJ+jkKSDMfLPaTdwPf7SNsdkzEiGhT2PtqYUwzSyyiMXPnik13mIUWrMbLD5IDqIacIBYri
Bw74vQZGNJwk+ArZmlkZGWw96nHF9+X+HZUJUHeZ1hPa9UptUI2OY4BULDkluK2qvPGXAvOGSnzO
rGd1uW3jkoyiuOJy2apJNweDd/uLOaOEDRgx1CrgVIEAVB0ajss8KpnAzeHN/GDRIhf4EEupiNxt
af3O7fWO05BV9YYPEG+uB5fkrydfhQAvt3kwFrN5PEtp3fQ8LQeBOo9gEDDgu3Mt/0Ro6upwFg0W
Uq8FEefUvg+EYf3HfTTUWNTj/If4W0cLmuH3Hdlz51PKLSW2o0+jPzjnapKPbHAO5WBH3wvszmH9
e7kVXV8rSsBKMMZ3qYmTKjPcd0Psdpjkpducnb46NjfA5vV7dd11aSANfzp1R4ZKoD/x9NXcK2JG
rFC2drt556QgZwOH6WGgoycL+VPHw8O62YqT11K0X6DQOEVORcSjguq/OJrfsa8H4QLgvk5E2fak
rdsm484G/hxpv2IvHQevW5Uw2LBv3ukOjoDcwHrWyCAy5CC3/xYpANyF4vQnWLr11JBLtzgnMt+m
LkaorTpZ7VcregN5AJ+pF7wmk6QT9yNKJvLEQ8zqqPTjpQdyW8/9J75LE416c7TPX7dg1F+0WIal
od6fGhiF2wQbmk9dIO9XAMdcm5BWSTQTePvGi4wkH5CSW400ao6bwbrXhx3sa8XufyRI9m3GZa+x
MclxIKJ/Vaa5v7k822xVrYn6oXULFsk2wDSaZVwzgYpPPZ/nQc4Lpvxw4eXw8rLqsQQB7c//vC+h
OpyKV0ll4ERGz7uZzwM17CUY02WHIHN+LyFQx1ZZ6wp0L+BXpfIokB2j2O8ez+VRyxpI7tgRPCkc
EioReJK++uNevdtX77kVRu8+zJA60iuvKexfzbC8B2JYIZaqtSwQAfcwMIc884tMRqXuj8fI43rD
TA3WbmQHZghBGGjYuljBZBQ+0/ylbvi+x++PFj4jOPAZ+LPUQ/MapupfCnBKyQnLGJt4GQLPvwkJ
mAFvpHTovR/7U5sCd9F3KdnQKp4xMtFEJv5cjzPjLFFtBv03AKomDcI68tXYXpr/dIiMwJ1lw4kK
CtNDmITsg+WBTa97QA/jwSfvXsRmWeZRknmYsttC/vA4Lk69MgMOJ4EW2z8FhcmxZTFGqOQm9ekO
obqz021IZBJyZqoWZiktlGRYJs//CB5bAdG5PGLItG/creAbRNWIdiI4Eu/kIrYZ9L4FBV3YXSSA
yiyhZ7WO2bPZwntGe5KLp+w0IvRX5Swm1CbGUAUCRnh29o+eEHxsqb9zd0GMl/wGdI4F34byOm/u
49ubo9Cufw7LvBX/LueKoePo2BFCAOfqGF8EVhNZ61Ct/I3myL3v4wE9LqukvDIwN2+7wDhwd+lC
qvlTs7UdtoMgSMZQ8YcekmmtugnmdMB8H9X3EhC9vdOIjk5A4yvEfBC3FEOT0hnOVpc9dtoyVMxG
dYNYOf8ZhwijV+AYEeAkkOk8J8muFkFmRhuUzesKd+v/Shg+1JX4einuF/alUTJP6+QWS5ZRzQu0
VMeL/o2L6niY5A33lsJTpEvtm6LVAN3xDcyjfxEUniperRbKMKl/AIr7o3keN5e8THx2yKj1azT9
2j49iB58iYvb7gAvw3w3HHxwJu3aflTQfplSJ2aNMgFjbdKRMPOapO3H7588OcUcyNLPBj76eIcp
tQObKeS8T9l+NgWrNTJ09TWtV/GYiwI6k9HPDfSvNH33phz53Ypqu9GK623icNy8I9Y9u9MwzdK5
OhRWSUoM3dWIdnjSpcU3Af5K+aEsnNxaw/BTtrBUN0DAneRBm7aIZencg+WdQYFQalMgmuOJmngL
F7TC2VY8PmI+x3NYaLRbuReRCS4caOkjLDzjX9a8RokUvLeyAwg8PzKeqZPJbyXV5FyZ/Ew+8VrB
qlFR2JGRQ9sT6RjFhXTodNspVwl2c5a3j1l6KxarVSK2ife09FGnnKbXJlu7wgcFdXxf064Qm1CN
5KLOMRcRRhWPBUu9FUYbeYFIocpdzK6USPgifmTW8V7Xd0QTtg6S54WZGpPM4pQSqa5v9STGa7Oj
tOqnQe1Ah4gMm8PyxWzfxQiU76/TndHBIo1yT3mPmKSaHQH4UIhTkVUrLfVXaXKsClfxFCnQdbWK
rUMDZKl+PAlMhCKTRVf/W4WTQiCzsAnKppj8FXgy4FB3slOG1l+RSCheUyGtotyKa72ef+fGLMJN
XomaRk1x/+sxd/CFYrzxa42cTYYN3KHBc9QidDT2t5r2AJGgaJAYp6sms9zo1p+NDHD6HzJzNqv8
ycdALk6mUjBMjd1YYRbsI5RBd+y0/ytBWZpX5ZqwF77Lmr8I5Vzc9YmbYbCFpChxvdunUNJc8lMv
6rcMfNC6GQplJG7PiJiILQKMgyKJkgOe3kbkbGJVxay0a7er4NA4UTYU616gnKfwFoXNW9C6kWjG
EW07Jkxgfh9pWR1MNmbzdxUqfkB5yjne5wwlp6WbRmLKinyrwHWp0YLkgNmNhmcMoIkCFkiYB2aW
WLql1HHnBn6N69qUu+NAPRwMLvDCaaDc7Y9AW9pTnN+jJcI0JKiQh5BUFZWmGW1YvNuJhTGlUbo4
KdpqbBptZftx3MdUhRjdVC7psf0rO+sKjwgSIMclwgoiidQDmy4EZh7CcetaEg4P3/ND0wCo6VuO
ZLoZ+SqVsZgQaUpFWZlDRW736PWdO7rxgcUsWeTkpMtzfik07yoLSWRmbjTQjQAGWvf0d9iyu9pu
vcdo1D95yEhGNL/jQkhC6yRP2bHqbN+ZTvia6lPnX1/gD+Q3n4dgOeewuNFDDkTgDTYTTFELvY3n
FQz2TjjT3cKz2tLEddSVl0b57Gzp9DDKYFxEZ/Sa2r76qbogPh3IbGIMobbE3sv6g1ucyaoqFPeP
PObf0Hccp6us9ZUkeQ8unAT6690VnU4QX1hj3/IhIW743X/9zzDL5w2TZrnxKUsSqI1He+7TWohP
rs6BdcqLzucoZ61JkepfSigv3VuTFPSkmK2LarV+skNAmQXbhz69pwF+OhaYpJ4v4b5VLnLha2TL
9136nveKhuqGKNxvXWU1U3CpZ0hQZwXufC8FPez5iNVuuv7ejKzhTalMo7IhMn1lQcLoSRRZAZX/
PyXHOiKBGyEF1DBKT6N1E1C1/tbDFTSO9PMY/3i/NqJZIIfY3F9mbJV0lVbl0OEjGRyqmrY8BU/b
IiwqvLG3JNCwcXAxHB+5MkHtJWPdJJCrcs8nVADAgt5TiEbE0opWK6xDuxyNduFvogCb7wZcBIXq
lTbH7hdfYu8DfYlTgw/YG/+B8dz1BGSgb8joncVSsUN0D/E9yca/9k798QEw+ZFlxjDUxwpyL1pj
gr/zwQX+nYGQeS2YLWLwBOwoiomaOMCopoPwUspLbRLQUkSI7WXToV3KS6dkv9+0dGdh06KZIcVe
R/z1SokAyoFhycWd8BLqHGvUxWUBxQ8puUf4yrpqWzCToUEMA4vSoxmI5SWhQfsYSNf0uUbS8tFf
HG95pc/UUjNifdE3xKIv/HYPT47YqyTKlf1aAhaVOftOpVb96xvuzOBC27Btd7Ob81YCLVGYv5Ii
I2cORwa0ybC663W8ET5wGymrC6jwUQrjT3MQx+wfK+P5drGXNY96nOgAJ5Yw0npjv7K616bmXd5i
Amdk41ug4+/NP3AwQT/JUcRrvi2Q994H0Y6Tt4Aov3BcljteKIAmwWlaFcwbzBsuhMIStUEUyskG
+zBpIvulPUebp8nnmy3UNzWr0ZUszY3utsUvXjrBI4ugCEuTb4WGCcIlGyJxGslzcnmehBkuYttm
vMxp1N5GPrDqujPrq2EnY2ovXfANPgsORzMJHPEvL7s+CJ6mONJWm8NSChQ06fC7BwQFaNNxZxFU
76MgFCixNJldO51ClEvAXDR/EttcBV7vHbWDzwnLRBvq+3FZm1paR9Fv+Q2GszwYKujmB975FjjJ
DPZZXpH6GcaZlfXcNndPOUxRGaCTG0m4YQJioxBCZEqbpTmTSl9zkONwQiXhrz0kMysSpYGa4+K5
eITIXFzuiKfCho3WQeHUXEFRW1g6wAacvqih10PXi1TQZPgSp7z3iGx5AcImZeJzGG/CvM5V6Ay1
HszjZXByt1gxFOsG7qEo0d06jGTgNihozOF8qYoDz5bWZPj6G7b98P1eATsWZLUUmaBIUGs1+byP
9eTeaNAxUbb3f+vo9EinujK8aFTAE042aIHE1GDlBojulTEsp9X+QZZo6Dba/8Mwyy47RVvCPzah
H/uNZVeg3DwmaMAy32LA/FNwIBh9X48aSH7oAaypUbjaE8fRQf04eOuov3JdywlBanzOn9Il8QUt
ECYqjWBJy9yzunehhDnj4mnaTuEATlPYDxT7rimL0bhWc7OUx+2VaoGVYm5yHHtCXTfjmIvwB16R
yUPFd0zz/WHobOmxm2B+QTqcFMaUFgG/QmZAbfuekCFZC9V/Tqx1+fexxhOY80Wv8J9hjjpfXpXc
qMAIw1fS7rFka5TRVy2faspuubJWSSMph5OX+h45KcYTVTxcMjgolqtOLgZddKotbCW1h7zYPx0q
m4rhq/stKqvYDev9LP2nLfbg6eN0elBS7wlgR8ujstpeA6tGJfF4V4CpY+spH34akTL4cCFvYh71
oaqh9DxNoz8SpjysUPvq9ncckuKPdgssTVfI1HpBsvM8LUEm/Sv2ZhnRHkOqu5rOfLrj2F+63vUN
AQ0WTfJV9MCpFeF43uFqmoEU1MStrbxwZ3dnAWXQG+BOotnj6/Xx18C0xHpEn2NG0kbugiuvSHcN
9BZabNFEgNVZ57jbcEKDDiWb4W/IenL4wiGddFR930wUQJ6m3z9zfD8bk1GAhylYq1Yh0jAdq4EA
6/Xy9Tp/gfqAqZhz9vSePKiZtgxmSG/4MJmuKP7rjwbaOTM1eQ7CkCIdGSZC7oBwS3T8iHAcviJK
erPLzCxMHb3uEy7Dx9YUdwMfuosfVTjNsLQdazC1HAGXjSi0ENMls7978aDthU+JFi1XQFkQlo+r
hjftTwWumf/H4GImuhLcQd0fgy3bGH75ypgBgI0nlFxO/tFuiBwQIZZahZ8QtVX2BjSr35jDQ6TU
Zadao3vDr44PIeSR5eiMnDEXW6kUuvq1V2OSFZB45PmNma+JsHoWhbgZbSeJkGoWdm4A7eqMNiR0
v+TOJuZxLGPftQsnPvlT/NGXYx8Aew0Zhtf3HSpOqaoVSCErl5uZXLku9Rre50bpOUYNc2eERKYT
XAxs//pYwAPvrLt0kVezpEgnMWQg/nNiE1sozhLjehP2gy9jH20Us5CaIYdKDChcc+b8/YJifSol
OhQ4MxxplTUJ14uZOCul0wiLLMoL5aISgAmpCjQ44yqWT4RiFyp/OgxOGgZs83iMNPQPGFCaD6Tt
pCkrsM3yBb1zt+eZlwdrVnx6R79P5f9Wz97ifJQO28nqiYKowP8EKpsUZc3Cf9KOyn+mNlFjT7/Q
nFBvALm9ei1iGZaYClxebH+YejLJJ+gD0AV5gqVniIE3XSeT1+ZiGj00w3d0uNjuOsubi3NykdCk
rgi2G1VDqEkRVLSjWANsyRkKAL8ymb8a7zDs37TuipN883ioKz3IO+nMDAomyz7189eKCoGH2ody
RXEsDSsYpUyMd8s25hwh9tFGctYVT7CDG0kNeluOOI3TWuY3aC2S2L4ZNE2bpEIijFndnVQVPYdN
e+TC0gHeNqEiaBfx205knzJJiAFDqYy5E3V14FTzGjU3f4KPZ6sXMW0Cz0ZiPb4QvGFXZSAoBPZe
OxsRvuMPRL7D3x6wGM6zYSozwOdAxxworUbeYw4QauITgLn4BsiXt8DPBg63Tgjtj/GpOmPy7g/L
w4kOLkNxYvqsduPUgI0NYqZR7v7NG+liv3kqmfnuHaEm4njzuPI9PVEXb70B7BpnPTe4PjoNOf43
tlRh4wzSNn8EbUclKcl1NI6M3fgXN2E+LrXoPZMGWfl+wUMGY+HOrcvpGPIuEP3Y5JOumnasFSv6
bHkeSjdE4OgVnbcynD3yH/MGFzQsg0imtXsqaBTPlj5LpaVdaCSq0H0iCBNhsfuhAVnr99xMCaGQ
e1o72r/MJRHrRE8jCBySs6bjBLgdJlF2Dzk9NppzdHUnsKwxmE6y1L2PkTQeco/dD09H/zLyTrkS
jQjLmFphTul1JbNp+KYvjvjBZrnRhVVH8YnzOi+jWIszP7Idf31HgLga+elNjyRzw1LGC4IMGYmF
9sK9kpvUhP9Nkkes6Sp6syKr7nKW9TYbfYqeGityiCN4Bk2RgUUvCuDm4tPQ6ogZ/mJYhUsbVbPS
kV7N7Xto2lECDljJpu0jjD8z3F8aY6ckFLrCi250yo2NLiTY9U5Vc+5aG/jm67htofgTjo3gW6M7
h41TIpMEQz9HVN6XPQyHH49HsbptiiPl9APh/nNtgZivORCeHH+GfM8ygssJOYgZznGUDg74g5GE
8Uzzmo0b15/LTNcoHWlQWEHe1DE6z4lk6KpDee4w4VSBsZnlVxsr8aYljlGEfl94A/SXZxm/I5ca
FGLr2HX0zRpiFxItp0yb23l9vd2H84uUdFJEQaWjxBqI3CmS4IvlsJtn3jsBfEz/EtsQM1aPaGq+
74+Cglyjhf2ERfkgEqK/4UNdzKVaWvrehYIzBNrAVavmnxcwzUpJT7iImHm1vMrKMqkT4WH6mNKQ
R1lYDYPZdvk6/ABTOG70Lor+MnjXSpz+J+EZCayZYJOEVoevjUN6tVM00bDTcz+Nv1FnhwoudgDV
lkIAYpz+wH+9eORFIGtrfwJDNn48IXMYCc5jevxUI0pBxzNNXqxRkocFTM0d8KAFhL9VVXqx9Ryk
//uFDDiUwRnaB2Y0D0mQcck7PCPQSPOpwxsjWCYxfguUJPHDRGQYVjuyE1Yqt+uUl/gLeJq7UEGu
HoBgxOCHO06G5ol23T/DqB5PpslG3Ou7IPiAyj4vwtMBqWgnG1mK80DL+9qjcB23BkV4zz1L+0cR
q6IyaKZdE3UHT2xcCpVSHH2CoFkitR8fyEQz6FAgaiDfjmDLwK+gjWivjHGjVS7cb0u2Eoww3YCz
9JabBQC3xiqJ1vVBp3w3Dz/9MrRSOKRj4/ehHfU1/FqxG3x6wFlWDjY6MIDADZJYPnViOkgS7uP5
EW2i1OVWhTb/dlHmc2mDSgLcry+GciTTTkfIkR/2BwmiXHI3B+KlutvVDM/TaX+piu3b4xnXbUsF
F8i9KG76+R//jPSZUyPpwQEuIkSPzBajW6KXdH6ttxcl6pYQLd+G6rjcLQPxFoek8nZJY+ieqzfb
gK3VLY2Badb/M7cYeIKtfoUSHJnCS5ZtKlkiNlgIkc+/PyjfyKmZM9zzbOw75OrdSV+h6DukzRHd
Zf35kQ4xnsliiCaE1vxktCOPx1rcR7GPcW/qG/0DksBrrQ67IrJDjhvXEHYhBYakqc9rUHHiDPCX
w74kL+8+w1Q0mi2h0soKmrXWvdue5wdTYmqYexlBObmaDhuApyiO95uEPdrkHNnawKzexYRZWsrI
KjU0Wn556vNMNCCqq850EeQXQLJ49qNeAb5/ssEr6/dfBR/IMKcvSbgXP8DUmUPii30I/nEk2vrh
JzHqFTLeN11apdjaodGd11Chpbxa2LwrX+4NS6g4xDqSpBCHLtK/Y95zyq5mgUUDX+rzo4pVvAUk
yx1WX9u9HUdX0JBMUXX8yNGP8wzWnZe1NQPgqUAlRXRqKDzzEtwXaqQxfoa+s1l7cETmJlchjOpq
JY3Fke84uQfWoCoUKlZqCLf3b9bS2vcxG9AsKkFgPJsVyqrgsBwG1qKceQKEGYJuYWn7rxi2daFz
ssI+GFgrUWMwLvaKdWt9KGfhU2uEMKNsT0uQzzC54ptVROOxE+KxjnA5zkktbKtiI9BqPTpH7zX0
NJl/omI1wvMscna0CuXhuEq/PGE0txO/npkmLYzbK/vwwYtUYnmQKmzdBSqvT/mngeDVTw3LNpMI
5lVSzGhkY3No0D3TzX+UGycqWEPuSbxkVy9UWnNLstaVPlis52HfxbI4m7xbzx+R+uq9QN5ucjEL
OHECy//u0BR2r4rg7TNwK5WpIygg8tgP61QeOEOURE1s62MWuYXPqkljzOgwfSTvZDlP8wwl1tl0
0985WItI1LGdvmRA82K1Z+8v2mypJ/OS7YDirQ+pdPsNqyCm9ZNnuNKUwI9zRfwxmwHV68oGQhJM
bRYJtoJV5IpwiA1euzHDUC8hj3MyUG7B3v0rXB0le/owI61J9qA/MrW+Et/Ul5XixE5+hO+3NXrS
H2Hmn51IZQqwRcLTW6RpdJpx9FLhUFlwEG7ax5IY7CEl7/aeT7uTtq4m6JXanA3ISgzeXAWsVVbX
ZxbCJ/cDXehroyVh3HCfu+TJO+rpzWGTNofQTIMjISSXrf2VNcikJXK2tFBgU10fzro7AsAzxBD4
jATkFyQmwhLXmwJbWO433tM4zJOwnPnJ1nspip9vGPikMKn8NQpgdX5CCc3HZV4/6q37F8HjszVP
G/v9Xw3BEa+gA6stpXMBhljmVxQ2V0hnk2Ie2wfpKZZ9nA5W8GVXFssWz06Z66j2U6vN2yV7wqyW
4dWQ/+/aWXxjiljNN5LHsgOu0WVPY6Yl3F8Y+yZOFFuLOrLrZ0yUj5jH9iC22M2OAuUxg6wUrmOe
pgI+vhXuYwAJWkVKvh/pr2b/kRN7+HWAyOmEPgDmFEvWISd7OJo9gRK4/h0h/ztb8aS28cHW9/KE
e7KKkSTW/TdMp+n21joFTqEl/j+lfAaZMM3XEX95lLcKICJksvAjEZ96PYIEpQxWxJLz6S4ROueE
MkIa5dw6BZmJrC37sC4PMGt+RCCQk5b3hSGHRrh7RAQL4sgpPprbvyHiIN3kERWXhqShqEHFTx6S
nkmkZpyX2BALSZf24HSKzsAQedgJOXlY7fV0RvX6Z8+BjX4gLE6LpS40fLMUJ5dd4+Fy3ZKNqzFg
KgxcIEY4/WM/qxKvnlWxiDekA6jylLJo5aQoI92Fqf3tK6wu9xQJkwZxjbyCbrMy3gXnL9e6wwX6
dvlHOgkyVdReb4sYn7qXhe3gK0/jPstu7pUXkqCp9XOV/rQ2pgirCECHL8NSHC+6cO/Infv9Npcj
m8lgn213y7JPwOHiPsD+cUslUgl0l+kW8Q6ciwMd96fXon8rdIEtH3Wk5jg5KndRmG9R1X2X64Rm
roYmWjenMYawY1np4xyiY2UagtPz8CGna5zZi1ogmrnjL/DSDctFhPlLwqSKQvLASSkxWAoIG0W8
lb+FgTR04Q/XHeCzegfjJojLifdeWwwDZhHrPjtYfv8BOb16F+gI1cAV01Fyc8g4iKsZVt25QYth
H/2JK4rds6rGaxvcyEv8PbWnodgAmJtgdrCKtgVViDnVZd4SLE4X4ZrIsHBw2GgUbdNYMODBtxIl
jCozuBojRSqWbwwvn6AMwWILUCYxsXZjl9mJ38CBudKZUcQ2R/TuTTRp8VQ/W9UimDKhiv55JySf
JRkbDKaJa/AtAFOSbESOYJueREhvQn7Agz6OqXvKGCojjljbLcEMDce0wOJa3oPZaSGKfMu6jN7/
mvPzOK8ipWILss/oNTGK3WzxcKm69CdmDwCWB3QG9s8xN1Av05Mc9sKLvIndxb3JkuJ6rqz9NOAT
q8nwWpYUkqg1wOxOsGkBKHKRVM3oyqCQiJN0kESDWoD4jk6GpAnOTLYrKoX2h9mk9ex9opfCOMRe
Fbgz3GRYX1gERbPhQVkxjMLbUP1AG3CrWbcmf6e7hVStEY++r02KvlKeSMbtjrVBjk4zoz1frr+o
DeU9uEcBRGAfLFxRZmFuB5rtdPf3rAgEMNUzQp7LQF3yzfr4hHGlTdu2eW9rdbJYYNCkOCxQJgBR
XFOvSo1EYo6TL5ku1MdCsQhr0geOVXeRmXkYLvVHWzrhkLyISIBfwiqZG3B1s9YdPdhCedwdf9La
RYjB9oPPe5AH5NQL81+oUiFeygBLZvdQ3hYC4Ycp+yoNwP/kGC9/3D8MfHxIfszAZMRPj5ZC0uPy
WtNl1WivDYafsMbon6tPEMH58FBsAw6pxym3RHTC4t0LaRLbZkt6h+loJdca07UyY8Gm2ng6Oqlg
/bpjQHULgmOsqyyZqyov4vUJIa2kVmrLOdpAkhmvwQOTFnoYnwbVK3gPeaoaL83Dsglg6crAiveJ
HzC7xvS9DCRCfKSbar79FzudbLVr/uvXovJPETEXrQRV6eGlIvRSK7I6F4HKsUWE7V3Mqler40i7
GU0snxMbyOAhaEyqZCDdh3EjkG8uPXvF4rsNrrzTFCGhUkY0/SZ7Ar+9770fUQtUj6GT1KZxT8BB
Uz1LUr9LFb3t3ZLqnLDVez/e9ndy/leuZVyTJhiz37R4TL8ZwEsNWyJ8oWB/Asgx874S8n3v+Vtn
d+SUdSA+IYJTUXeErL5Ffk0q/ZfUO3ksj954xjZq70EXG8W6ai7vcdQkiz/yQPkfU4LvpfFSrkZd
i545eurd2NEx3Zin9YnCOeI5qrxjFa/7ehZ41+cSwpO/McECU6RF6SpJkPsdylDDzkAogDnxrRRy
zMZ/cfWF2JHvKnnI/jD4eWnGUsufXmXHD3Qvjugttv4g00HluG87cRE0e/uORdCC3tnKhaH0aM5F
tb2OOx0ZmRzC/hg8UlXhirKAHNUL6fdMFFNhWXUaZEXJRLdVj97KepctaVRG0YZaczyGwNokdEcW
lS/NSoK6TMeDRgIcMKI3wtEnlkj+G6yOg+Q8y7ZEzpPYL3gd9udxKDw4PmnpaJsujZQIr86ECx0d
/9QevubBsfogvJ/U21i4CtTxrCdU/FykCIOwdXbM6IxReXJ+u9YPH38rqEp1RwR5xbJ5kCVOHq0j
LgN79UnBuhPWCzf4K5/A1zVhWzt58VQSzghJFgXk2ISjX9SMfemfyUBm2SkNB++SuGN0Mpc+Y9e/
rpPTPlAszLnZjCa47/sWWHF9RJYIjn72Fsd910opX1n8Owy+Kpm5feTjN0l08JWPnU0k2qxiIt7Y
7TddiStuoEijrUnJBBdzdf44mvuJ04t+MgE2+aGZQBdxb41OjY6nKAXvSm8rdSM7zbSqoGvu7RBT
rzx0K1wSB9ys/VfDdERqPcNfBatNUd01jurobRYmg33eLhLo5MWvOkgzUXBkA26M9AEhs7aFDS+o
7agsiQRaXAKBgW4rCbcprxZDdd0CToPJkHvxEvPBE5LCrVi828WBhhgomd7QW9Y3FMDWHHGLq0J/
OQC4u1t0hHUQgsvgllwlt+MuNBxXnn2v1iJuFHXDm2rmotGaUmKhX1Pt/SfyFi7lNKXnIge+G2BH
h6L9o//uBwrVkO78zJGmEPxPmfZV9ce9o2HUTxSJOhlr4zPBduM5eQlU52AROyI39Yg2cZqfuWzf
3XHXqipuckUvH6NHeVoypidp7sDmF5Pgf9gaGpvuTjE9QtAoPjo0X+CW/5UVZorWEi8H/3Jd3Kjs
1DjMuOo7MuDKLVyfnO5JlHzv7FfA+OdpqneLB9VEL0phD/3mrKI6NwZdMNJKBa5mCrzoYeuUUcSn
nia32qO70ffdF4Feajf4aHjHqLnhbI4UZ+XY/mC4aBQXW6bOpsNRlrDJPFjP9xLGY1ItoMbXe0+E
UOpPInFJOXgYmmufXBee/4oF7XkeHpr2xDaA+J/wEUPWv9RnSeRtsYrmR34mejmzyLet61qFcFXu
avSVx3rJPYFGiTXUAmAjBK54gKRmSr1zcwWWYjQv4qjFZ3nQdvwEKyoX65h+lXjKzUP5YC/WHo8I
cE1mSKcOFc4ZivbGEY7ggnp3gnAebOXSEADcSt3B0jZyfL0gLFu3kRtalDUip0D7BN68wnJy6nAS
WnkavAN3OVT1Mo26cJQzeTeBBZCMTVaGt8v/00NEOU1PKeIlJG+fPHm06Z6O2pOda85eB7PvtYgm
0DmJ8VZF8WJ4vDFPOZeyg21YeJPBUlZTZAAFbSNbzPd3GvDIc+qy/zepRSfj6uDProPahiVDuOPA
XPqFm4VKKH/NTdTKZOSXId+VPffmbvt/LDSiz0ycOj0W+T+Q+SRh5+MiAzvRwL/5mX8VuQrFFjPX
axuMpv8xwLyU9VI49JT4DObJgfRbqZYIwDsEZXJuOGgxAY3IM4vucLbJBPLai1OuyaBaXX45aeB+
HI7xbwFVj6cmkUpbRCoLtcqd6Wl1yd8YQj5/uD4TvwRjhtdAtJbG6xT7ILoMTPwP9+IWWYMBtByc
bsyrcUbqm6qm17Gn/lqRCkDvKVPIahMrReHxH1XGNf7gqnIYMliOtweQiafOwKit4yqKBZKutM4m
wXcKvFORPsGKrnzEUpY/vk2KwYnU+tBmlyBNXfCZL+meHMEOwKyClKBW9N5JKpwdjGCCltE4G2lK
3PEzj7duAY7uwS3rQtx0COd24tNMtNJ3EF3KL9WT3jFDpx0PzhaloX/+oqOmKvznbNkjM0MDTgGX
oZxpx2er+uiuCNArf3MTGTanyGlSsEcNn7u6xWnh97NVK/OeEnPcG1En+zBqP2SOr13e/+1qJAIN
Glq9aqMXaU+/kv9noLP/T9NXLsNlbJ2MlIkke4FlUYN7HSS6e02GK6PRTn4zCxkkVtXqId3FucP4
YOKs02xssZPhl+A6WYZRQcDmjdb2tR8s9qrEvIy0fr6g7WKMRPmn3ksgmxBS92YPwQ8mCjK+55jV
lpLmKzc+uVPFRfAxaqJOefwzqOQ0zPYsAHPMz8YTFJQMzHBABZISy+nReZgv+PxoYaw1kBr3P4aL
aXhxY0ZkjQhplb/0cZFtHx/fC49HYbcdX/wV5uAPU21OS+l/V0HdktH9fSdX7FM8m3LQUPKCIs5e
WJotHpDiq3ghHivik1bmYoLp4KlVUeI4XpTapZ61JbeARNN0NBhofpxVne07B4geDU2xclUlrtR8
Mat2X1gLwctxokBv0Hl5nBF8WlJhMvKMTwkiyjjJ/d3WllpH3uBFGgVfSQ3F8UOX77ST3xBPMboy
YLc9Ri+AM7ZBzMTz2ZSq9NQZaFZjaZ3nHeLHuxmbqnYdAD4FyDIaH5umgPf3SFqbVp6c8jttWtJI
KA8apDr6KYHhe3lz+CwOR/5oElY1WOnhs+WGC8Hq6IbYmaFrOGTjoh0ez2ZiWT3QIeqDHqtpBivP
jyVIchE5/8cUBwLsdePssnZKv2Rss+TvjVJ+TbVgb57KSee3z0ptqWJn/uZ63TaSD/n/5oNFyfdp
kxfdh46SezQ0NpZAhyyi8YydgZTsZ+74xUCWtiIEtltJrLM7vBCtk8IuYXdl5ywYdklEGKHbKEbj
8uEjOE8Rps/lHEKh5jDHk7GBP6JV1SuEi7gfGTr8m3QGleCdfCq32eqiYyxr4RWjWTf9aDG1J3Ln
2rSLSsSMbJ+0sMsROjLXBNgpgdwdtLnJiz5a2/X767unVcPcuO60OPYFzPdwwpTcuqI9HbIYAa2U
4bF67vNk5Mm5q9vVHLKWPrnLzk8k+XMMGR4uOb+rpWfNjxwZZZm/G5o0g5cXlrTYPPl60TNK1Shb
cR3ag6sLrgla7F51kACKaUGc91RWU8RRf71NSX1AL0WRYXCTT7aauUjAUzZGLlqWeV3TEljCxk28
Ni9nyZRCHACSvjl/eXxeEPH50eKCHLHDKFd2hNQgag7xiFPOD1OWLLTMy21XcKAYCuZm5mvvJ4gK
3G7/a00PLBNkThRjL3ARkPK3yXcwPelgA1ZGAd81JZVS45xe7RBcuepFBKCKDHQeusaQb8VR8JB+
IZlLhDXgZZggMRG++vSS2LNaJWZ7nTbNd3mT9mTjR5SWzzlhPotcHIWWMsBdkLSalCpzkILT/MHE
qQNNW/7nS6mrr4if9SkEeZaNWVtYPUvLBEtey6lJXSFyEX2mpaHN2QGoyhbvnnFxz2NV2eIaYFs3
9r93h7KHxOHGMq9r4CH9iaJFzEMov4SLX9NDdx8AOlr82V25bqzCmJbz8/xxxZYRHGtna5tlH5DD
OHlY8sLYkm97QdM3npc7DBLPmh8giJEXZRpNi4dzDVru8uifKPHuYYvo7vRy/QGx3xd45+tKE4yS
FyoInn7m3tk49e2a1s7SZHbYclcmzOMl2hVqiKo0hTcTlEDX1rimm68F3ZnJtN87AEiiGb7PtijM
xqtH53aH+3I0g5Q+JIq/FSNOL6C2eiLG7MKUpAEeAZ1NyfrUltfaDBqA8CS1enta3ctrGHr3iI/N
bMlak0ZKA2l3xUr6dS5KoUcJsC43XJnqV86uffZGjjnqRHRA2eOsdpNKJY9pOKsX3s1l+R4LO9Y+
JJ5kilBcIkJfOJ354WcIKGM2TY57mS5dofOGJcNePG3Ve9mvh1yfzSekVcf/EMG7ITdmznzj2qEE
ssIbMBTtDMzRMf6pENFdo0osPnMWqkqh2/Gni+GI/wo7/1FUAwsv2px3SxWbJj8aOioHZlxgl6PJ
O+ZDnEmn2g9Bhy2hNAdzy7VMHo5QEPWn+83qx8AA1WicKUD33BJmtGm3povNon9H2Vom5m000rM+
LlBmdEeIUUZgqHwJuQR5KrR0ROCmNnQtpCjzmcNrYDaFEpP98TAb98SXB5KLTHx0sXOjM8tfce91
pKXuxpnJhu32noUyYZikB2ycB4/caxu30YdsQ2nmaPxWxUnR4wKe+g8no2avbNlsswnwkM54N/K5
D6oODH0yZZIjG/s2WmHlZOliccsB0lVYcqIw3Ep2bFlXSwA7sSRI2p7tUgxC1FHgqjqfw7Y2aoGX
l0bdY3wZKdbKRhZ4S4HopMSwdHbcCfboBRBC4sOtR1Qe61Edddoe9zES36AwyZuNMcy/ioEe5A+h
6pR63tZehcs51T1FTkeufQmfJKkrify0puJ5+CW4jIK5j6f0Is5Yt3Wqus2CY2HJypwBXfm5xjDp
TnFyAG/gIo1DJC20EFETrysMfMnCMYjgHUsDDLPUCF7Ri3hm5NnnqFkBh8UBleEMTuXaf1k94Cq0
wfnnUhBLXa8h4nZG1nDvk0123xlIjj/xMRDAXPVLmNYRhQ37ohTmm/wg5cuU6SlR/UYOox6ZV6RS
+smu+ZkS8VAQegG9FLXtDBaz71oy67M/C2YXARMSDkfOS6HikdlCSmdkApn4vTvXYXylb4xZYaaS
3bxW070hNstQYOgc2MON01PGJt0P7AggVXCZAoZ2XWR2X2ZEeHHBm/9KSMJ9iCxqs6bMKiV5Q2xj
2S1PnLE5/4eAM/6aCGX1J84XznobeGlb0FgP8VG+dMn5SsuU9M4KV1UybjOld3uVx00LWpFv7Z1S
E/TnjKWV5/k5CuptAJ5LlDnOUOL4dDrN/ND8FeIHSou0lcwN7jzWPDRGe0vyIUZgB72A6c1XMWYk
/4aB38D1ein3hfGuwKbEbxt6xdGfLg7vKtThBTZLLZ+T2pjGN9pO6phyFo0ETkMKgA7oHUB5AFWK
jm4txdH2RWM1uVTcFkxkMCHURSW7nZ701ftLKC1WNK02frSF2PBWaoCzXi5qtelPqYhcQH75ybZK
9nfIlMlilsjLwUSbcaE8HsTHJySPOTJDcgesfLOkKo3nnW7ZYYG2kc4vZBBakwMOq08KgfjS4iIl
PMtkE6MUGUFyeEypEv/EL7DnsxgGZOkAKhFIy+TLS8CtpbenF00NIYnGJ5oXC8ARbTSVP6VavkeU
Bs4qlmjQnJPW1d0zgqTMCqo/s87rFf9l7u56H7LeTpvmHXQkXjz+lcRHBUl012ihzQMtEEZQbh8O
CrcEtSfj/qUnvbwMSwKgAxkvdAkA5M3fYjWiqx2qVhYh49iCHaNGlNEMCfc8W4dw2QYZW2UJSjAr
y5HW+aExrqptr9nZFMFRfXvStUpa7xo6VKumy4WtETZUWCqUPfrUgxlDdfU9hWwgCuWeNWMcf7/b
/efzWUJjyxyBdF5Y7nDHXMN5O7dZZ5ocQ4qIbqYGNYPkxwrzfbROLDzl789l+ZIGupy1Nfcfc5UM
UdvVqRRRZkgH3MsRTHICYBTmFDZdWalK0BYPgGdhtmCqCt02Dp7UuQZLSbJNkdjPMSqjBfP+T+cG
GEJqLaqE8+X8uPcUIhjHiM1RxNFr6gkpZD7A6iD+J3fJcFnF1GlayrKWMOocgUxQ3DgacUBIhjQs
gVNHhk6oHsWRnhG7MHPScP9o/LLXjdm/aonRj180tfzpBinEKGsEFW/w1bXyzzpGgytYAYutbmzU
54W6l6HcdzARNF7hyMPfYpNECAIY8+kba9gR/zv8C65gwa4LXzQ6BUl/TH6F5zZqkaOG0suu4kja
5mprrn9aJf/wCagl9Du4y8h2CLsPlz6iS/t3K9ftGVt8q5bPhWMHZAW33Q1/pJu0KO/bxHIXwOHw
CFjKqLFFJDFz/tnoNdO3NO5snIhnCQUtP1kD/BPzeMYylG/Qqoq5mQxRmafv/e0NGGfVAxRVOMEz
2cPXc3urcvgWpo9RRaTi+UnXJ1GkDjFRq7B01RWOHB4SWpSekPsd/CjJOQFg5SZyBMCn55rvNsVJ
AVNJuUyfnH6Kllp4Fp2PL0OITVqez0u0udPgPHIGlwnDeRg9c77q/kXCy/nUOCeeipn05FUyDnUA
uV6s0VXK4TrnEZpr5UkVqyiXuxtcm8ZOOEhZ2BYzVv5mvPgsy9x41EmUlpJRFzsXuFMuqw1oCOZP
DMp2Lkc2thaaRYBokIyxnDsoSxRNuVEZtBNDDK8GHoD7SVOCEWRTxXKLoz7ahSwglpNbBeDvJnAl
74WV1xmbHmdejK9n+dmx/R/RRb8/UM0g5yZ9onDHZaddI7YLrnB/Qf9rJj/6DQf/KXyBb5ZMhgY3
2OvoZLb+/wRTFaocAb2e42Ny8EkKTqegtXDL3CFDyP+soXKxdKiZVzg3U7CVvrF4vxx7lHLyWJ13
KDkL3QEtbkRMI7ifdRuGNT13jgadPTFhY3vCesJyEOUSeimg/bRcsxUe21SzzhH8PcVte2rxYk+w
htFz6RaQofnZvgVr2BkWbFOKuARbWQYI7aZD/6bAyV5tLWAO0RB76R7Z+uUOK7QMYQhAaI5elFRp
oNCNgvVM1PBTs1PbC1VdZbm/gBpbzBvoZi013WX4+tLBePtwDaFTfOTgzFIHnaJZ4POgFVj/Ibd9
jSKTOj0cmyVxSv0e/7tHuDEyY46vi6scRHAlq9l1P6I5JxFnhU6OS8g0FssSVFE4lVxgfQRP9QNd
ayeXUGKIVfC6VM7u276vNEmoku+bUrhH7lvmLZYrd0qbGi8QRd+hSDHeLhp7Bwlhla2wHhqnCoR2
LP437az2fiWGsLPUjycIWygPGTEVpxwybne/aqfAoc2OdnnesUr2Nu91/VVt/nAANA1WT8FnpRMG
hsmni1S8BDhI96TLaZm0T/zVNc6/XNAQNG/i5a1mzE6xNuNJBozfUDWemejswCtf+IWlArqudf+K
X9EKvC1HELgv79JimZwFRgCbtFMtqkmNVj2W68WfdzM/x1XLOKH0xaQIjjs25KE1PUVJ/SVmyuvQ
M9cXRLlp2XAYIMb1AQgTMDJ+VH7En4ILQBjxa9pJrGN/lU/eVsiTWJQUQjoVm/TyCzy/dpmNzYqQ
s4buICKISeTW7qaGwS/3kgqgfZM4V3yXwtPkGsxxtb2Y0V+7PUf6TYg/xi2/8YDoPp2OmnEn0sYJ
YLXVuFybosyETpuYKVA/XLJuk9A+CrGfEFLFpN9Mc18RUp1eqgbOy7T3kx1+jqwEOdfGhE/My8ap
pWi2MwSVreSLvAnkQwYsdCbk4B8YlFOiQXdmu3228q0egJ0CkZR1Sx47MNuNUSQBZ8uXBHOxHKfd
BAD+u5+gGTqBk7rYI6+CI0h1zrWtV6g5yhbFXxadmTgWJzgb/pV0ZIW77wxqFeapvPj0q0Aur8cP
f0rM+auQSkUdB1Q2yFaXHwHiIolSfk5JIHsw09YFxU+zlMBfaEd8j50ifhdXtVelul9mnc4zahfG
j1eBhz5vnlUdoCeOfCD58zVf+0w68GFvahf62ScnVRGbxMVfnmrhS0R473Us7N/6LUzhmo5OPqnc
Ibn0ipElaMl1hzLs4XpV+oM0fyxuJNY0cZ/l0A6OXBZ7Ft7SAE4yd//89SU1IbzGptGkK3aMnFZ2
ASoBA3Z1qT0MPynf++Hfpn1jfDZTcZzLLwODQbXLv/ox0+6IejKZ2vl/i9/grt14qr7jf34hB+U7
wkIqGOyMOwwmKOWeTqfq21iEo5Tv5DD+1ebbXe87lKrBOi0QYj2KnfKIqjwpLNBKH1QZ4doAGzWk
UhhaC5jnmlk++ziWRaG6QErRJXkqzuQ9z5QPMhRFT+ukbeTMfCY55Iq47Apu9tu1UGIxOQBoAaqC
iVr/H2r1Oo4RvB4xWRXK1ny9Bg3t1h3aiy19LTLGP77gF/H+rYBfFQZuvIgYejjDaijRfKq03ATh
VD0VNPXjydGTva6fCVXX/59fIui1FvuD10BxiGWUEXss4SVHWcqaMw8FIwCxUbrnu4dGqyd7O4NF
XKQNy4koK0H4GGwiEvhmIThPb+z5tbP9wpGDq31Rz7gD1/uH33qNEKyyjFKTPOoIPDqzpp3CnJK0
wRO//shPN7b4vA86H0KU9Uoz3qa97lA71YH+/3Tp1RQ4H4qAl+NlovL+41e1Wsh3UuUvNIOE7q/h
G+5qotGMmQ0ZshDlfoVd0u1iEv9lBig1FSMJjFWWJMMExBvXpRw8dl5C+DiSDIJqokvxPF8GItrn
3rD8HCu/62rTuDyveqXZo9OvdlDyy39zFstprifpEOjuDcrMHChaeMiKpD5M6re88fBrnM5DvoGr
K5dyCRDexNegBqf4mjIfcOibkDLDMipKZTzpAhZovWMhCRJvVosomEVO6cUus8T/g6qxkAkbLtPi
eAymVdZLdGdAzG/rpHHpRT5Qip7ggYtxZfHrW6iHSRbFtQ2kWuJ/oOUska7h/L6UBOX3WzX1Dy1+
DREAj5aQWUJyYkpa7SoGeeKA8C4jsCO0IMaMEJTuorMGPrcaipVb68wotBemJIsd0HOV4JDrL0Vu
jzZDxzmzRrAhfmhj5YttHj2nQlKj6CrYPDrU0Xt+gniD66qveLzVD2zipZCVNVQs8g2PJ93aZbvi
cKy2ZwTFbz+dnFAPuo5NAsTEtAHho+s7P0Z2txj7iPGsEEySuMhwCoPtp/HHG0I7QEjG5F74uega
aePfGpK+vs/RXBKvmqBT4yLf8PmTebvDUgI8v1G1rTY7owB3BTSlIT8TCtCCMBeDOtPVy4DHpj1h
0K0PrNmcu1qCBiLwxQLZeJMN/tssNQky9fCerzCJedCFY2Dcv8wVwYfykAsPIpwM2kecauSqPsUs
oITHx2pt3cnCbFztc5S22t/Io2RUkqk1e5kx5QzfsPkwMDk4erVpi8R5QYUlwsXQ488pB2ib7HpN
Ao9h7Wca6Ykotl+6z8haP8WMLcUJUiBDWCbydSdHibSUn+XnsPluldumDAlGNUJDG8iFRrynq9/p
UxK9aKqtYC/MgVRda57muEfDRAC6vxuB1ZPKIkjpYvS0/Z+db4Sjt29shell76aMbBzwSK8RpNFH
/Zb3r8l0IXUTjMk9/Od2RDdpw/JvFLr71QsMAmeqPVteIVYZzZ4dcHOCzGvdPCR0KEBPqrBXkPAl
OZbiJ3hlbsKuXynY3Ub0syOP8EbjbERI6yVZOjvuHEBAXFev8dT8caYOxLdYtlprkLopc36Yb6SC
qucJBVBeqrBSkG3riw3zplBrlIs03HoVYiq/kpS1rIVl+67jt+AYvNr8I8uYdeaIVc7fGxwDztsP
BLCxVrodK7gjGcBf9f6eQ8Qq2SBSne4EqybOqKOkAalEtzRzB3BWYI1Y7/fnGiLEWsjqW0Tfy2wW
Zp5Ho9Vsh8VpwjnyEzjLrfWxfPTAqZL2l2LPhPeHkFGXsI5Toc5s7P8LufeeH0gsT6KZGmExrLWS
hi+tNL/auLMTOTRAo077ebHNSDHxTocCVsyyI+9iIxnIE55isvUlGY4H3tW0a6bZJWEaePB7GKiE
P4i+IS3/pXzjqYRFoR5CSw+5hb1j+OXa9D/5rO5yp0okxJeADnPrFk8xJHgVDcfHfKiPwhnBPcOT
//qn4bsUr2WsFuYywwYabxdmlJiwmTY194M7PBnVWKVXFvI4maZL+nzL6GXfiX1ACgV1MyTLJVhl
rSUPZs/ZsNcKH9Vcp51Co4XZTrlvQ9Q4zyrbVqm+y+bIR+Z6LzQJLywLs3pUL3dWTioz2foncRB+
ZRqoc2iml0Xn+XLnPXud8Rw5SAXoaW6RPMmF5fbwtCspv6T+FJoC8HHj4eiED0mCl7/U5/EwGCjP
Pi+sdpQnes8v6DZHvxJKrzKkRZ4jCqQfBHbwQ/y2kgnD6ZcbmgSvDiFTXuQyC0smDzOtGPfjlL5p
sM2Z7BNJCQ7mNuDCYItgF1dVT3avWo8bewwIFx+r0Qa0YLhjiSZTENrGtkIGYmkCOzZYWARVg0rr
CraWdhcGlLCsTvGSy59mpg1H3O66Asw5UWnDMmehAJH3EPgRGeaEVvA7Us22XeSKhe5SePpNTd3K
PoI24gbMOzkMeU0Gf5wbNXowSoJ1GN7yIhFDFAU+8B9yH7x1hnup3RhSti5TnNYVZQ47QzcYdE5r
3y5Zvc+fG8eiInPcQphjnAyLNGy9fVxoW54mWctyAWOFx/6ngRaj+p8kfxsLqUBkZENwXD49Pxx+
iCLFeiy3keC+JnzGI6Q2vnTbD493CqCYZxv8Es0B0fr3MAjyWyy60AI6PHBT/KN42q67shwqLVe0
VDBIUYd06DA35saFfPmQfoNhmPaxPeACu5QShdi/Pju7oR5bFch2cRuWSb+TrH4NG54hFUa5h6OR
P4clILF2INlHnuCg7D8JnuKQ99Mq8Nn9Fi9ns87AdDsuUZcmOWtaVWxywRuLer7Mf1phYrVqo/mm
CMQx+VQekdxgfjWFOzBB6y5YOCdonvxcd5MBuf2PlRFRMl/1TdxohTu7B4szkdsx3hqNH5n8x6Sc
wSlRAN+bu+Q3oo1X2qMSY3vyqjeVa0yNC0UCEIPJ3nKHA4hBcp0FJeHa5W9dxVNbOpDbL5lZtzEa
r/qin3QzhT/hZROLJYOvGXYuf+zfHUuemg469jkMg0OIPlth8whsl67lJQC9noDL+w4Zh1hveMj5
ycFzGRw7gpDVnjzVlR/lpVeCWtpTH+EbggliaocJk48WNUrpIUWqwnXg6d9XmuHv3RKK7orwRt/e
lptnN5ELf8nJY3f6TVhVFIRY0MmuO23XKbaNYwdzUuw0IAJ87VqjH7sEUPlUPKaQ6AOSi1IbkfSo
eKq1dvW5Wv2fS9JYt/cKNT6Gfe8lG8Ap68imzZ8BgAyIBWJ4YmDw54M4bv4NaLSUgxG5eUzYcOcK
cVH+S3J8YgNa6OokA17BHQu1YoeHzbKOQDxBAmQ8WiqbuNCZD/DlOTklcMBn8WmQmB80fz/hBjMQ
/uDqqBpfN0HcNCWifY5SNfulWBYNkjQotAqkjocPRw2q2JNjC0JNNpRiY2WxuGPE6/nKrVBw9K3G
XlFnvoI8IW9osp9IbVzczWXypBHIlnnsYO8BrOETtimxiUoibLZuYJBm+03glgIzAW86vx23JRvp
FRisRoESxfDUYtjLx+8cEWN26uyR5+H/mx/hsUX7fP73HRuqOO6h/LFh4/chcigfZFZPCnAJgR/a
tR8reCr2C3WmKyPUv+P3b6Xt5ob+KJ7kmM+y9TQvNwW7Qww6faE/wLGG5c/m3GWskWymnEl7qIgy
saX4su5Y/f8JXSTl8d9TIR+ixrlieY6+3JXggb52YvgUtvDDFiamk6+OX6SP9ITYM9SQxfUCAHax
1cUCpqj2MfDWjNJtsIWoyoxWV1OSZu9TlHXFJ0DdeLzM1nn97oicseC0b0aMvW5vY0Cv+JPxGjv1
gxmpPBuB89ZCaoT9XpWP3lC7S4NVPpltWkDjzZo8CH/rqtor7/9E/L/FWsLlg6v2yOBQWJoHgzCu
8HZmrxF5Apf7gtsfH0PJhHViDj3NjW0ccXUW77jgFZJP3eJCh+UV5OMFjA5zpzsrJoyet+xL1AlT
aUDVTHZGRGxt066QPCLx4RXM/34AugdtYsjqNzvvbdU7ahlS6yTMMV7xSk+Qo9lSWUwuyLtvyHLI
+mdHLvdQLLP13h+p4k3xAGsXOV7H4z4+x2JJ3jWGMK7UuMwxls8oRgysZmP0gqLC58UdvtHYKOGi
XUOyfp3jizwkZGKTIcTu7UmyqwCZtnsG3TxDfcIERR6El8kkAgbVGmr768nGVT6s162o6UQqJpsY
opWSjNoX0Ty7g/h9tayBIDIUWPcwQODwFcdN9WOWdUgOsKH7TT4urQUFA3ND9Eg9qLyqW1v60Hg9
Lmc5Uab4IcdfYqAz/dpPYUmEfVAako2iEMYMBcflatdb6JsZQ1rwYpzkXA4T1vy5ChsxxUcKvKrB
GS/gCjCblr/I9GAY8V8hySkXbyn3/hrLKKZNoKIfI96RPgWvT/viH3AwpdPjiSYSNFhVG4o7+3sm
e9kOQafs9uv1NLK//nJcZgD5FfwmEwbXwEghuDI1haxkpicU9t8CdMWejALCTnLPt/H62vRHF1OV
rUSgTxNmSgjzZNRbuWOyhKGbqcUI+t12hzlj311IwkTUzoZC7+m7WZj2UgZElEO6bBfsGQ72i43s
tCUG1mySu+ILlqPBRB7XU6XnInIcpqhn6lIsd3Pd3sAob4XkbMOzJEZ9QH909LoxFJC0dbvp+NJO
JoBD9IMkVS1ekT6kEiLdlHxJCNJM3OOi11gCkhfj2IxlYGyuuaic/pGl7vJMiA7porRYxTy7tf8P
kMI6f7gJmwmRwAg8rB6Fi7Kyel97hH9O24FLP9uoun3xujWOSVMegLYYTh1rXSi7uc96PiZYTRoY
xnn+LITC138awqwGZ7wwQx+JhhQjeeYrrwI1sNkIv/L5Qdfjz+BZudpaXztD77kNMjyuVCCfMwSq
yKBSxk0dqL3BRMPoZBJ98E2+ylJQY7j8arxIVfXQr8ukhai9p2f6K0PRFDJkbP+OSgT7FfoxSOkj
oyEg+gR7mRI+TEfiKBmlmEZQVTNIsKNGeBwat4D3TBAbctNNZde4G5Ww6vqqdxzA3LixldrFtetK
/6zhmvBaqP5VIR0M/r7kcZxb4ZaIvhEw8ie7c+4xfwIElU/YIJ2XvgiHGfV+u8k+sVao5wAz2FTj
VSM/w4Xf8qzaPvCYvdVHD6GT0Ru5mSx4LoglG7mx+OfMb7J9ly12OvbZiUGlaZcTPpQ1FZ8zEbbH
T/yrqHrXCkbbbTi5uXn+zx7sT6YgEOZbBq+ppg0Mv3QzjUFsbVhmrOTm+hTDzC2MPTbsDrywpKRC
JSmtqJRd1nUHfXJOGzymUQNBOkgJaq3boWiMxTcVB88zLGhFQFBI7JWCSLC1xcvG49DqGLZNfDEv
HbRYSElJZlzwD1oucj9g1jhayssydHSrIdX3vU9iNHhmrji/smL/6QR9LFaAGI684IWXhqqaF49Q
xeZiz0hPG0FbE0gmOFw/3FZfg1+eQvekexSup7118YvXkD5Uapq+wNahm+8km5Inw4ZdYqSJ17sq
3TsUCwt4YscKa1IxzL4f1lxkeSr4hAK+u9BnKAb/TEsNEz6ryJ+7n9mJSl9UbjCcxKNUppAeRJhN
yDZg6COiqlDA4ZyOVlmD7XT2yg37cekllCTZjvhyrRAdv1hMi/unPgapjiCELYITOF0mGKiySzUQ
9RfcnWdAk/k9zxSiDy0TMcs9PeXWlya30YLeLoNvj6mRcP1jZAYbKlbXHyMSaLkuIWxAt32dGnNM
T+KTIBgh4kThp7AnM7UmYZ0sinl7Fn69IL5SywI0bu+fg/K3QuP4DgWVTZ6divl+4JumDMePVf/X
gyQrPhjZeK2n0aX/VEX8NS0E/WrzUjBlEW1pUNZnpQureh2nCw9lPs5OX/yo4hTXwxjOlOvZ9MW9
g5e62foZZtC5y3g+4OnY8H0rGG9FF7r3hxqITfwSyd3kOKgpfaawTQ4GwY099Ape/JPG6b0MitNv
ymDiRHwSx9WkLI1MWKrLuISxiGvFY5cWRIuxVtbct5pp6xTgEPFt6JJWuNsiu1rPt5iy5rW+kcXQ
jW3ok5Kh0nV5Wm7fdmzNBiw2tepbTGjzlvJJDXtO4JFVBwpciqn1hIL/pH2WfXh7nTBrDZFzZl2A
uhesQ7lSaJjh7Z5zYNS8nmKoWWm/hkeDkOBmmwiO3ZyjwGfEuQjWmycS/8ZvfFv1rwVhcaVekeYr
USz6Fbg98UffJd4jpyli2hzGrF/IqTshRCoS9Dy/ZLUpjWs9ErQ862OQZz3/P7VXKIsPvaTwUFPK
0d7WEIL6F6AV75aeqh897HFmygKvKLBguh2c7gI7zhM4yOa7r4bhi3BuUpA1N7pJHDZliw6C2eNZ
Otm0ZCNfS5Dl4MCAeHN5/sx+1H98IE/as6+x1ji8unNGDUhMFzGfqHlNqQfBqCjcsA4w0KjdwzPH
vbbFeig9SUCxQlsy7GsJH3tGg8lk/jYT1n3EqmzEG5k43tmpcq5+rL3hYHcDitLVLvU12EAn+e7r
zzcoCWuq72uWaQxMh7VtlDLraHVwmoZSuHS+fuiL3R1vABrjwAdgxZ/luRPKhaOZOmdycy4QtuB1
T/0oU8HAT3mY5hSxl8OPNfr85Kmi4JJTQ0/fila0f0cAN9nb6s3R4OIq6UzbK8v17+HGQyE61X+P
lbAWYM9KkTWTbpOS33UrmgMP7ejuM5GOIcy8QTpP+geW9Jix4WHD3BKam0LCST+B8n48jvMXLmxR
Qtfc1buT93TPDRIBOnPRW84F9ClezVc2xEua/IE5ZoaScKqabYXKiNF+Nf8syWdTTMMeQkKwi74A
aSQrrsmDss0WvzhjA3S1RbT8MQqK9P/JrEnovNm7heP+Bg5NNo2AuSt2Nl8uAn7BZCS68/Xtq5JY
Jxc+scfj2V5Z6SNUgsfAcQz2MulzYgLz+3QGm0/6ztL4gfanR7N+dVMGyM7DLbjkEvh9oT9OpIpa
zXbqJVe47qAlvQaUj/jyp3xLOLnFz2faCZMOKBlSAa2XMAe3qeHAthaqwk9vZFO4cQG6I+HbHbkf
uelcwbwe7iZHx5BwPNaf+jI8QulYpnY99DlhtFeiDDmj0Ws3xsNq4YOmzXexkTKHBfpnPrUz/HXS
jhxw2C2uQDJM2HgRnevu50sIoOnrhicgqNFiOyOrrBXx0neLJ6RPZ0R0qqvbnoWLOLRufNw8ucr0
G5krvmp9aSJSD3CZsUYpoQ7181m/JEPVSbBZqLDQd+i8ZD+UkDO621SUOnRhUov4X01c4+xUM6lg
5rJ9mnlbBgv68Rckn8RPcDX6kWMCwg3wvmk3MJ2sdcnV7ZlI3R7nx7iiXi3SR2h5tI+322KwopOm
3ORwNe1Mfs2LowtxlodZzwfhQEqNcuIP989Seeax2DZXORMD4wYTxGiUt+jgPdLkXX/znchLzpdj
o0tdoxvF/hzHdObejaibZaEsIdj48rQ4uwnaJteIMLR8m9GT2wkd8jqSUeSrCTcHBv+xwOxfkP1o
LRmLgyzLUDSj2afA3Stpufu3EsYxTHYVusKI62y/N7iVeSN+8pNApQrwKfYKeguxO2fC48wAhtw5
Uz9J6xLyBY/mt7288vrnxFTD9tPyIw4bvxzWFIvrAEDHdGDbAjOmacZBsfzpV+33Zf1EHRGXtYvK
K5KSQ/3xIIrGY1OThn4jvSA1KyL9x0IXBlM/TPeHa4Klc++gE0/+W+U2wmAMTh4bpyY/koPP2lm2
+V814oYDZ+L3sh52tarNVMbBuEA8OshhZWIonVNM4QU9dlgpv3GwMFq9kdroLLEMzr7nUb664u4Y
wMa02+NeTe4ImnuIvsUubf6QAW1aawCnuBknHwmFzuiC5DAEWsi6fwJvy4FtodSZqDlk9AVFozgy
dqdd/dl0pvbYZhXYAi4mbw3aIJSd4Di9puCeeKRYcpcnaGzHHGdIC4c0GSKAHY2xmCZM4TyUV4Fa
D1I40vQpzFVQUv7WCKWk2zMi/f8aQ1Ttj1D+TM57vl2m/+leacOodzSYb4LM0HZ2DSjCxVNc5x2c
mg77iYIfyiNx8njleCSVNYrvOYCLGH+z1CviNLK+dSDqhtjXlJ2ZCp4FpR/vJ0sOB6Su/pgCKGEi
Y0S067JvX24sJUWT/abd8HZ+0QuuO3r39OQaKDWImNWD71nsmmt9XxxgnTTC3ZEqJbv7z3MtuJH1
WQyTeci1kUT2nU81n/0xSqRDql1wcoUG9TqgHmm4+y0gsJ9v+vIHyQ26aYn5o3wbud33uoRmh67O
8cclv09OCUZRngtgiPEu8qgJQehxLk41lWuUvFd8x3ujRGGFhIYT4kdKzTfWTPOReYuYSfzu/Wfc
p4g+VB5KrhnPCwTyGb+SP+DI9crx8nwDwtkRgFZ2oI3PT679n34YpDTCzxw26UUBwdO8vRZC9/hg
rDOMb4DoYPVG2cPLTIUafF3/xNJ+bOBZhgfyqZ+CvZjdVaLSkMkUuR+uknvjkDTSkhbluVIyunVa
sXDMwPU9rEm6Gfjk6zcvwcZ1jCnzZTYCHZLY08IfM0R1/1qeOSvaeAJRQ7qJdWQMGo98Awz2taCI
jLpVkF8bek/CrUpSz7gsQ4OipAojHTOMzlOo7gTE5bHHFkpmSCxJKxgzdQiEE6H56XM5WBbnCFZp
dQeyheMOsD7m04h5NWdOLMWSlXTYsuee1Ll7Ol9SJ3TLcEQegrDeC5IlygvVOjsHcKwhS8/5ZIzJ
fPEJGBxGfV9wqWzJ9TpsxlsA4bhPG8m5kSeFZPi6BcgcyL5svWJ0GBQ2EgG4pehbsTZzUbm8UyJQ
4k5g0a9msjj0gdxmIRDJ+LeltFyaU3iZDLEXIa2XVYC7qrnuG6pe1J9wK5AXJ3JtyaD82qSVbdor
dD1gwO9YYRLk5mlTUs6LZqbQI1QMs54w2HcCdTBaNMeYiRB+7zOL4LScIfP30FcXhxHT/Wl/cI3g
ZgqJqAE/vSYhbAKQFpOzRHr0Vk+igLnvtN8CBL2+qOb5JRkEgKf29FpeOUcQqQe1/TZ9NHU6CYEq
HGlR7DaHhGAHPdqqqGXC8bLWd1Q/3RQjwknruqrZkzbo5AjpV6hoWP4eXclQYjHzkcZk68uFw4hH
xqYhSGNeNGt0+qVxBdwE2mXCKGtrzOw7QltYBM1ThKfUDj8xBrasMdpcpqNgYoSXZbgF+S3CdMgQ
d9Jqgx6oTMk5DNRM1N5Ffivs0Zu+4he/4n1MwAOt2byDSnkL6HMJPIr6ZyqCcRrCjrSYb8b/FlfV
W8fIZ6uaAGW6y/qvBph6LWfpEIkpABnoz2kK794A5x7cMosEjR2zlwq2QfmVxP42CbqP3Y7TqCM8
MrDSYERxwPJoUTIiCcsJvtOIUTnXMVCqbg5lEC+CZSCYWkqAOkGkpexPtBJsW20a7+lfwztXMQ+C
d1jKqfi7sD3I8W0wiii0/Z5cpicLXkuLVy3u9V3X56GtaIeEPuSfQhN6haV1bRMSJTwH1EFj3U36
uiP1n7lGzS3swzmgLqVUk16n6r5RyrmaXwE59nM//xfq97UWYpzNTIkXP3NYYFQ7UoFmMTpbeRLU
C9NGNf9L5K9csPDGMiDmH4uWwaCIN+pCPQe8qQ0m8VisV+QgoA0qTfbru23nlKAdJwnQk4kGNgiJ
wDILN9/kgWECVLFpQsET9VwuOPF33kDO/PME8F0h/bZzXTPxPND/5oEiJu30oeWBJpzobGk5rpYr
iBVC6JJObVSTSRcYuAiWqrM/25Pi60xIv441w8z4/jS4ypLxs/j1aC7LLsCu9zDqmGn1+VuzT/PD
1JGjPLQr+FA/KfYIslUQeUV/mv9IRbzcqG/eHWudi/anmoP+x1ZgSIwmuP+XZ9TpevLoWURRPUvY
qhlcbol6zkMI5AJwDk/+i4FSENwuruyrJ+YawfuMTW63dmAeeHGISfJJjQFhNjHthcAqGzMlleou
kyCgBbpOgduF5Ee4af/uC7Y1/PUcZrv6d+YPGlcvKNtJmwPXBiHhqxpftpvNC5FR7tF6AAuNCGOV
PjmyZPlkLxW3KKoRMEPKSduItfFWTUXPNjdL2L5QMe9zGPIQ0/SDrYRYMKr3MaXAcK59yTd4pfCj
pLfOyIKvVuUEDfuhw0f43zG5afw5JHnLGZEjYzT0poz0wJHe5N23U8+9vxuxFdDhlJovNr9GYsyP
kLMR0K73pfedyDfItwP8j/bT8y4tb9OV0DRsFXHQ6VbBMzHdf+rgt17CpUfAZP65dwHHjczhk7Ta
719e354P8NIXL3rPvCz1NQeBViU+9luDS897Jw29KCC51/m7YGeoSEDscIl3NAJOBnNOnU9oW3LU
JkSiuT2kNZccG31FcchUppYtT1ujHDKgVNWP1V4IQpUXrkQ98hnfRd4x67ncVPhb44kKAPwyTho8
PE17iKSY9qqpLfxFd9N0JnEvIerVugl1krIc3KrTJKsxx7fb9KIvfPDh7bg7chXSVIasH047bHJw
tDwMRL4JdXVriyvhEtVbh7tsrJwZaMhFrSHZBf4RWee0Fct3Mo0OnVVfHm55o9NWb8USz+Rdx5zU
6ECJZmnLAmGRbR9QHkrdsgH/vGb9e8Ov4FCctZT/l2YEby/n7ceYKOLJkLxAjoYM7LTcggsWuOus
93g/bfAImM0bwt2goBKC0Lz1o37++WU5GAkk5B057TQku4wUXWfNhAjB+JfZ8XE+l4ii9J2VQBUI
Cg0tYIlcPuOwt6aDshNK1T1xQl5ONU9uad1Zkq0wnQqDQyayuabNvMAJQxeebJfmmGGk+ePQ/C3l
dHufHsNfGhozx9G4VjGRSI2R9vwjDi3TUjxadujoxini67IU/RpDdnGUm8bRyEuU9L1+jjmmm1oC
FNfox45hynEppplKqu/rgwcicaeqr6EntSwQSng+fumNlFK4F9U1uOiWyOJeuYhiv5C9IYehmiZb
4ELAk4os5mVZOb0ZvyvXq+5NDZ0OwH3yuYhXb5M82art1Oo4Jw3iEH3h8HH7ADkqpAxDgHqQbgr6
2dCe2ZwKa8rKa0xG0cLOCNvQsOL0tl42aXujqv1QPoJ/prRyigaEq/DAsiZCH2q3NDvNvCTvukBA
fZ+dPypGHOkOLkxrfmmQfochhfAncBXk+0jE+HT0SEA7I2tTX+0W9bD8B0b8unvkWlPJ8P071QW+
dVG41+Hbgqa/aYAXnrqPQEo86izwfIxcHfrT8wziE2Ef/u1syZ0lUZwAdMDaeQIjfOS7/7RSRSsb
+Ggb4hFpDenjQVboeZ/5FESsphwQ3LH49ZsSa3gEBb58eNwMsWkB3TANEs4dp8foAgbmwCCqSEhn
lSymsPYOIB7yJqDKdEMxrloOXkYC+QUbkzyMs4uVheXgkLymMo2B9t56l6t3mHnavIhClOCVOc2U
VMXqyRGWVxYBRLqS1PvA593rZAJcKD9kko9BL4XYWuyi030Rd+5Qk2ISchw2qGbrZ7jKuE+WASE9
lseEvGvOpT+EQXGWoO7x6JAbTVtjyyFCJCvMAU9UKcVxf/jzCkCVzDZdyP1uMSB5Eff3qmY0FGLb
AES6f9O+E0RuqMQp3+rK17LT6V/NoLmvDChUpca+hAv7zgr/JH8sXr83aCIK9NtA4LaysJ32eNNd
WzvYWFnD2dKtoX8Rka5lihDV2udcXSBlo8uuVGgkP88f2PKBcMRVkaRKGOiwQJwwANhtLr5XoJqc
b1hbn4gqwTjUppSDMY7nOZaTnirQ/qIAiuNyrk5Ru+MNhyDx1phmPnwag5eN54AujthaMHnvMJls
UwhQFFxQYKVrEAOqE8czeEaQ9S7iNDeZrjy0Vxa6RGMZmqGBb8DYZuKh8zI9qqfwXopK5DBdZv11
mGCnnadLHbsLc4fLniCU2qpFlKCkMWhfNHjJgfKxbvp9bTlcfFVjZZpEzONNaYWP1qTOQ8/XsrHZ
LZdvgANI+9slM5Bxh77BKkIYZ9O04/suf8vFj/iAzCHPNf27xdlxyZbv38xrVKGM6lmoPMNBnsBZ
OVWn9vxEeBblAx/jgFQ4dmyxsE31mSPOYJphUesiQoE+1ht41Msz0SJrXt4kMXOf6dvfbdYnIdRz
EFf9GCRMF03Av/pA/WdW5ObctRn1wZj6kAQQUJhsFli4fZ9CtV/ZXSd5x0WNQmLjCmaRySMJGhPM
1tMxRU1P0w4zDxa5e5axlZBB1HjD5WJgFVINmwLW0T+rXlc5M6VlCa+1chy+cXq2iF2Pj4f4QBMd
3vRkr9wvNRUKreUGlp5/A/KhhVf60gBcdNNxF2c1K4Bhd4eWRvhgvi7CnsCnfDamEIsk8N60XQCc
FEh5CpT1FgjdrIzGru7NK8MpcZ9+a7TfK/2LcvE0Maa4nTvODxar+oI94gkI1//4Jru/uFzmc8XH
ov03D99cif8acvW0+4azVHm7upXlziOSSa8Ret8meV6N2sfgz8/QT9JjX1nYe3H7efCcnmUMpnUG
omx7nqZu2co1WFOgojx/aCCNLwbeNeboDKKT+j1koLQ+bu5dCEvBolXZXkMzxQRs4foCeZoCjeen
xiaHX0o+v+Nt/OkhmGnuh/DBZzoyi0573iJc/owVgb+9Sauh37trxTHovvN+S9LwikA3EIopVaq1
7DfJJDtlN7eq6TUBri7jLeUGOkW9yQMfg3r0oZrPUD9BuSRh3CD92xJCiwY1f2LVLtBmPM4GqRRW
2crYwJYIc3O+Ia+NGhXaWBb0294+G8ab3s1egHlr1/8Rto4gtMhJEgBVU0RTSaVuoWACrg+9DT+N
2ELn4LolKTRsQdzbiV2hKUCVmUo03f05I2TTckG8NDjHANo/l/QBU6PGxoIl5jgea2P9DfmWMu6Z
0G16S3+Zp3FeyQd8CMQDJT4LY0eu7yuBSfw3q1PEBBrNf/dVr+ZfiNHVg4SIF9mVl9xPim98YVRD
tJ/8W66O/a0oiwFXBKEvWMtzmR4zMMudONBoXfFojK7jUa29gpKrzXwAHlkUBjLNRnoK8vZ/2rCD
VDBmTV5rwa2QJMfw5NVVoBs4LTM5K6EDB+dI5A/JQ1yVpYr3aJ661fTH7F3kG47UsSIFp/RK/pRH
+zTwlqo4v47OIu5yPiLHmUYwK/ITDp/Z7+x69di6f95wqu3EW2VveYYpWZn7MJIGvhWm7sefMPcs
BRSjx11bpV1A5nd14oMHwR7Csn6Zz801tdz8l+64Rs0m3Tkj7YX/fk709BOnv/HY4tYPOGZbVqRY
+s8cCAa7r+KqOkt1hJ/02WoQ/8zZAeKQ3QP2+5S/HsL9ePLqN8CIW3UVBfn2gBr13Zob4EYMyN9l
6xrlv97AcZyPhl67tnEQLnYoTFZGYNDuJ8oau/tCjBdenfJtaDo6ryCnlWD0DM9wxGSpX6cKuizH
xnf6WNDEEwIVAHOG3Qw972zd1RekmQQioLi6cfXn7C99AMEdw3NNUvVa9UxqIPDfho89k07gAbC/
vmptdpXG5o4VPaQwYYE4YDn+wjNbSJ2LdbanXoJDH8plfbiDRQy6e3IgYAEnlAeWwUef/QABAecS
JdAoVCs1Nt56hYdDS9aQudcZe/ipESEioZVf33InUVhmgf0I76SR6wy7WFzVM7ubu2uUL/BJg2dc
ihnra7oHJVqja38qNXmaE62ab2W8xOpo8vha3MYfqIZtp+c6v+JRzfi4Esv0+SA3AGm0/xgQDsbl
h28YkP+5uh2Y+rIvgccxMXoIYfciIo3u3wwkb1xWXjfcuIexUqSOCWzjTQ0FT0ZtpPp5fAuju5uF
YnJXO6d+ftIY1QkdYNgSFP8C9hk9uf8vAdPWQ06zbQYFZcKvEpbHtpDCKtgeXMX/0cXJC3vVag4H
BbxcHePTqVpouaZiGPnTI0pImFGCD/WaJbY/30Km05LmZ7Jkyf1W/UhYAgO+FR31vH6CE2fax1PT
mqsPyuDKxtI8EzwCNkkUQF6sYgqoVQ09nh58oaWJtZMqzrC7I14RPtzSGQar5mMHEzIhEaiFqxKY
XWZgWdmpxezZKKfD867tbd9L4DghY/cP3rGfTa13CpkYESnIv6ievkqrxxRcErT2zEUBQkILenny
GJpnpTJpQDmNOuVuGo7k+nVJJ6lKkXf83IIDofAOT9+4cDepbrByzA+HA7gGh39F4u19RoNU1FBt
jKjv7XX1zMgWzsHTqiVnTdeaiuUo/3bgFQOab9NH34BctLzhDx1JTnr68elexxqcde7gm4z4TQaB
uXx+/ROfRiI15SWJbJb5rR1uSe8PQ/1NceqE/NNE/VvX4tNWpTFhqEQpHWc1EguTOKpeXzMEBObF
oWBlgJ3TlM81m+lB6MO0G5K0/53a+y54sqGZj3EOrcQB6+fQGOOC5TGy4/cNCyBHSoTha7kWyTPq
XKq539zTaEhh9WBTwA9bO5lMzZEeAosZ1edya0rI8m2H4mtTWYLWDPAjCj7JwpL1V0TdgsSi8MZA
HAKLzsiFxqwsLdEg+dj21d5EQcU3FWfLtTCLcsJHQMJmPU4UjTOsXu9enjxGtEiNFyAD80CocIwf
TkBsIuckWphjK1oK0xIWrHxUpWh2Tu54Hv7ktMlr9RBiuAwsBTSfb/ZxY81uF1ayehCX7cPTrRsS
GSLeMc3+coY24SzLzIL3H++qUlB+Oe2Mo1GEbcQoTPTiX2psFNM3U8TDM1Kioe5br/2cOaZa9WEv
k9pWPjNc+Z0/qyU4yLgTFNfZP5eGseXjXbVBASgf3SmUm1qf74+bsVIXJ8e8PCCNvA+1WaQBd1F0
CWmVS5IJf8qgNaQfr+CE0UGMjaJa2g43brFOABM3Ecla+sUNYY1NdScXqBUEVTDDFBGcMwkJ6onD
agwnHGhaAOYMhm7iFgWR9pBxmazrhshGp4pIT2UZEH6ZNh9o5hDAfGqpnjWDflMyv+Km8mXpu58z
z6V2/0PJktzN4YU15x79yw7LN+mmwUoK5/6edKcgOLHY8n160Mtvr5P0uKTUnLqaTLQNr+oaALxS
UbnXyg6xZTY4EeLCU2feKF8ir6s0Cxch2AeH4n5/0M7dmPm1IZMmu4wlCdVXFSXnzHFzZht1Gbd3
rdGcLlnbmyM5cjUFE2djmjMijcdwo8Dmmibi4sISAj/rH8HXsTtGZjDGjJHuSOepDQKSmtUREHDn
GkCHhN8EzFALjFaIox1nwXmnHV/rEeuccDL3exygFxXsvm5KUIlJU+MieTC1/JlBaIKUgwJMsuAP
zvnG1YEOyZbEiZqJJrCeCdlW1SmwR/MAqnYnFVUvipPGBTiB87RJ/KC+mfqVgES1uwE4oTeihvtk
BoacAeaW0CbEAKW5BQQ5YIPpwnVOM6OVXh13KyggXFBTXVUeUsUOrV26b95EaGxNTpbGntkTBBKV
/YRUUA6y+ijWl7uSEWOMNE4QiBET6XNe4+kjCh1MMYuly5zzsAJc0acrbg6ZOI91upr4pYdqhrwh
mZyQwv/0zCbQJApJ11qVrIpbeyrfLy1R+xRTBcL0JQiyRmJqdoqn7Wmdk/1LuQO49Kjcgjaygc1r
pfNYfKhuGOb1q+mBXmCmLUbmuAA4PHin5HMYBIm7Jdhpj4/iIKX8qY7DFTgVf5NWoH8RKho3SuQx
xGOnYHVdeThDb438mnsAYy7EupVPvduaEA5VNRgBq5w3LguAdk3ROvWqA4O8MxYoBYPe5T3phwah
UenrNT6JVN/n3/Y7dc5G3sC5NM5eKLlxsKyovXSh+x0Jztpr9fDIIjdSGd1MA+bLrE7O9lRJXnoL
IT8d/ph+uWtpHK6tvnZttPSLH7kpP1yntiVBx58H/kiD9YlEeKFmg6nIVfjFBEWS9KTb9knC/iwv
18XtVgTSdn6r94uC82ddKveLsNJoJCwfxnbNt5Z/jDjF1DQSEWZnfsQQgKADwtVJl+y8413AtaWd
+PXWoQyYdDA03ul6GVBMNIxeBPF/fMkFrytXnY3/kZyciqlXD4Xvj1k4lNzcMKxgKKDNGdAYhtp0
wzTmef72WCGWffhD1tcNBRw+xu19ZgstNQPCJZiOU1svp5GCfs/Gc+r/lL1h99c1giz/Cb0Tmv/B
0WtNrKC5t6EcAXpqUD2+CW3A8qTyYm6fjQmL+R4dPhX44uKfJKeQ43WyVsOSKHmkb7pnqz4Obizk
RHZCBl14UEfJQkS6rWJC2WFG90kkOJkI0mdI3VjG/yaP7Z27lxjZm8tz10gd2GXMc9Y2ompgdQzg
H7gjBfUU8bJ5DxATscMgNAw1e6WEV1kaetr0h9LMFo+M/UhzmPbJ69rXw4ainBPg74DC72TIH4sC
mbxGEQeXRWTSZWqnKnrm/68eP8gX2HUqo2nxg+IQorLSuyodjyqO2IADTWxu4LJjYKuwsn8HQWkk
tafGIEpB+IUG3i+mmDDEsqLQekoqhmRYzNhZlkX4zeHT4EX8qIfusqAPd2Yus7HEa4ddLom4e39I
PEs72FYnCmoBKfb0HdS5R7Zq6MsaMbwpmbndD1RHTeM/70sFl4uKNe0KXVqUsKJX5jdBlivxXvVJ
MkXa3wmBeC1CDqSuJbLJ058O8jIyFRo2v9c2l4hJOPA6EVd8H/oTY/0xA/gON/nsy/R93CA3K1Mv
UD5k0/1IjTej3au9k2FmLGBFZ2nu8mK1MLtFPngbmj/HkAGubwKNYPNd4WKmnU6cuC/MCV1dlSJm
hMAPHCkKqcUkUC0mDcrDsJH4UEZEEynDu2QLkm9uuDISIYRw66EJf+W++PQpq/bBrMbsIBU4wq++
BgEBO84ZT1fWtEbtZoZQz4T4NfGaHAvDnx7NQAnXvhqZ93l7djMWxENrZBMZPdHSdhLOIg5I0V+j
YMBshD/d1J5j5ANdlUHx0+y0UGVt04Kz2wq3StxKSxr+XLICCmHB2GTDfXzFo8hCGZTEbdtuXqlO
jtQxTaxnw3IpwCDmsTnGJX298Uekx07ryHwvakE6us8a5G2a9Jlk82A1pllg9oW5HEwyVLbXuJLi
0JUyZx5HWVbnNG/SHKIwNSNzdNTk60R/a3qUehHGqgTF5k8v2iXzFTdb6SYpR2/NbW3FIEu2GalH
WiTXaK6Sv7vg+DRNISvkfa7ZPMXt0sMqb2xQ8qyFakiHjj19Yj382pltDAI2K9EwV7qWOP+g9TvS
lbbzlu5BxQ3WVuH8N5n7GapdjE7WJ2ar/Lvv/SdTUx86cDBtfoJDHWE9vFNAz1LSgXeW3cwR9Aih
4EuxDmJWVDOodr016yN4XCqhgowJZ9ZaOv0J2dP6WZSKLYwdPacClT4A3ziU+EyqV9G2cIbF2K7+
9NNTP+t8WfAg79uVTM65V+PnanStsiBxf3G1spEmM0cI6s5gTGjXZUq1+l2//29sJ2oyVWWhqYSE
nB332qvogEO8j20KG/aZp2rPp2KSX06d0Na44QdJHwoFoCwIYpdgZa2c7v+tuSKJd9svh9TVGhiQ
MRqYSWCQytSqv0mhJ/asiYCocmZyxJ1MwSTSeq0j/9WdkX9epfbN+fQfsNLaap7PomScSP5Uiamg
NKFIn9FGkRqI+sEJhXspF/p9l0BcrXmjdeZTuYoxy08adruIm79M6DAhLWZNRBZw/OJqbfNlk0X7
kGVqJewYxFbAtr6YQkkzLPObmJxTQZPiOze68mFORKIoxKK8G4Be9+R3Rc4/sNRVKNNxiVVgjwwE
ArKEUjbpGV2YN0/vvHU6J8rohjyr0AT5+kkHluyxrHmoiILREWrYOmsFJU2EK1JZuHKeIiIrNsIJ
mgwAxYoRvDUrkW47877afRtTp0S6zHfYH3ONPbL+3xzab19CM4r1KnyHH6H4gptm49p6Ti/zuvxA
BjQbXnnvKwVuJXDRIC4CH2d204Ddwm0Mcvlnsnaf8/x6YRpOqXPzqQipV4/3gxXfpWn8SLSC+t9c
ZNYOLVGN//7alf4f8CP+OPjkvRofjz6YWx0ILt1D7m2CnpbbkX32XboE0oTq0GeuGjmAxLbINiP4
Fp8WzEIrOonZ9zOWnQVIclSJippb+FYuUhKsU5el/K12cDFrMuIvIO1TnXd3sGDXNbMRLUA1GQAE
p7JJ4f8KayOtFjEUVIEDr+swbgOL5Wc8X8FajMygYBGIHE13CYJYnuva4743ASC5cja653WGPbfk
b3B7FBJGUdO1sfUuGQ7Tda0oqvOcU6J/6o9StxZL3Iz4labvfFTSByLEOAmh9Ry32Ov0yduuxwQN
r5EoON4ZP1c8T2KNNpALjljnt+hwIqg5ztzK/5lQ7gYQ9x1wV8ivqApwBkVhaz9Tge1UBVfH4g+C
h9sR+wEJYhujI7QrgrDXHmPsCR2uUBIXgBedDmoK1HHsyWFXnlZpQ6G7y62BzQVpFjnvyO3ogvKi
OWYBaIsSL0q4swZUZUYN6gDIIrcQJpqd1eONg8MCe01o0F/p+2K2wdzDfdbrxVhZY7dv5ZFANLvK
CIzCzgwKmLWQVrkGsjXGywhidAXcCKGuhoSAFtKDIeWL2emDRrnnj/sAil1qIbzghz207EynLHN8
rjOZ1Sqn4QAuwECKJIz4CD5skV0HpKLqLYSjX4H60R5Cb/Hqozyt22rVu+/2Dkb66FR0WQcPBWCh
UYTg8TNMWID7aZNFlRFnvSFg3mom2FGpARNes1536Jlx3Wk13Tx0fEhMZfPbEkIw5+bSetDFdcIw
0/G8yh9tP9uLLD463ZbyiHtZNDa5lEXJEJ0r+IXhOABlGT0pLGTkTtrMgvigsqI0WlQUyn/Whyi0
12Rhrr5gyumkzGX3nG4SvcXV1R7tMOcZ2ldgnyUbX5A0+rAQWT3Yh1948ScfgzkVPKwIzXet+xLU
SGrEsGlVk7LY+2vw3ABPZ9ciUr8gY6UMvj8fbVmJR0HNvhMU4kvv4J1/kuKk45Fziw9yJEMdikY6
Yw3M8ysyUyN2fqQS6gGxU3qdImMnBcuk9mx0lEPO4nVizMCrCVZfHq1ZGeIjr2UTjQYS2dD31SlR
cajHKUoOBZ20FVeaLpbLkRglNdHPNGizuUf9e7MPggPk56b7FyFbPOrMpvxjHbiJLA6LYn7d/iOR
L8RZN7LtLb6Bc5qK5rs7foiyTRP81H/iSirZQLVOtaZ6wHIIqcfdCUKUAZfiMBm4mPrwFLXI+bN3
CER8huAkoo324WUvPIqNf6QYGt4nfsh1bs5IQ/a3PXOQocoRrnXfMUbgWFQYHZhwWEKzZ186S6CT
/Tg941TnLYywneEV5gqylYSHNfe6j2S5zaprt9u5iG6re3wEq2bRUhPFNSiVsF7OPQz6bzOCePZg
hi+raPqvd16xb3r/Ip7ijmuY2qJ8q9fO38XbSanBnSBVTu1t3Af3jyikPuntIIMEkHDHxwH7/+j4
mXYvr5wjGePHYckn3x5Hw8Ns+csTMS/F2X51eBEK9Iw0/0r8toyYcFcpqp4fVmpzu3Z7Hl4jiJ6+
uZKvkFBez7yXSB88K787e9Yhs6ChTGZ0UL+ivVZJXOUthFwbd/19Peb/heIRNwjf5hSYFE18mYZF
1uPcrF5ZGtuwiVCr63vFNIDFVagq6oXXc7oN0AZrNEdSsERX8jgdrnS1GhP1tZRP+iBJ7HKFclgo
7Yi84lwdA0NZpnIQUuXmo2nxmCr5H8zCYPaqi9hOH6Zb02gjNxr1Oew3qB70L3qnDJfMt+jZcsLA
4e/B6pA4TEocZP4DdpoRNg9rSvWz5zjtMC0T+q6zCsO9DvttJXuffsFCs0KEduTrd1r1FVr1dJWZ
WZ+xIwgR74MpT3Ufy2mqZl5H8awQlLfpBANihy84RmUOHeeozJIvd4FnI9PSOCATtBinu9xdPLQh
su38zVEe378Pd/d86TUt7J7kjkGDkAeMyuQkYXVLsP6d1q2UnB6R8LLk4xlbfv5VgmuIm9fcAXsx
KxT3XJJX66eHZ3373V/gbEhwC/DE7V6Ll53FTmC2H8ikpRyMkJf6ITsBLKNK5kUrzUbkVoEsBs4C
8LPCMFCZ2TD3YsdDNhFl+3AUI24SCQ1TN0fJRAQD8tYsBnqhVPec7nh1lyjf/c744nMYxDD6F9R/
gzN9O1XFi6QMgrUYRUlZZWNBh232pDguDtyJ0J8wF/cwgw79DWuapPKieZ0/K8hG3R9qy6YXU9y2
TUK2GWg8Snt3dTXz1la5pd7Pbr/dGfMpRjYIXDf59wO+yXHnrpmxLGpIQm6jSUhHN/RleRY0RlDv
t02DAwmq9yR9SWi/NaBJ2lE+JEjVt/u+518BWztZTCNxbZswhbUtMaS2//qBBDeTEb4h4i2Z1/ZC
CLBxGJS6t0QmKnj5N7ah6RS0ZXgJ4840likXSV73AsdfMd54T5aLyBuLE/DCK3yf6RMgZVwpLTBX
Rw4uPs5FoXq1HVVdNLGCb8EApCsiI0CHIGC4WSGoQLdb7sk0+bePZnK3i//Msavl/vc1ffr2OITe
qRwVOgOfB7AX3SihoGnhoRBz2yyzgsFdlmtAsTC5sBPgjQu0o2FOAJd6mMD0s5K8zWSfEqGVsPQR
zoDzd6o6lv4tBqRoF7CQaUXTGsjADek31Qd8keCkKEartU5rLSHq2bMPTTUR9vO1idng7sRe2CXE
4qNULABfhWRd9GKNZCEKY/jO6Jw4TY90MHWhpNfhkKcbb3WZC+1qbupfT70J6cyXi4RfSe5k0a6y
m6oKrr6pjBhePNo4HQdQtURP+0wpAuPd50Fock+I6gRcpGODZ3sHozZQmw+CT0sTnHkh7mK0jOKl
BwylKkrFQVzY9kp1CL6ctFtteuK+FQqaKxf/DIyw0F3Ba4Dd40dOjDFfc+6HxKlx9LpOw8PcXIDA
yzSxj0PtfDS1Hba4sD5443vG++nIfrRw7Vz5MCkUn/iB3ZlAHtJjFlROZtYmeGjoUsGNyRHZkd/v
0rH2xVeuZEneiRvQsJAk9C9AP5dnutEtFO//HtCrB+gWrdAuGIbpmmzZlRUO2sHRikl+rWywNxQL
FaWfhiCHLk4RayQ7j9YqHC4orlkgw08kr+5pE9mg8Ny3iuJMPvv1hcSFlXtPzTr1TnqhdYEBEA1r
rf/mf3u6qAMx/qPG5IsHQ+EZJmol/c2EVK6KLVRSALuka+b19c8n4j85/ZOGY98VzU7Bx3IuKD3t
1Jpghy83R/izwKD6qm7bZ1MuHJ9Hegn4FSxsyeoGF8k3EnHCMANClmCN9iss0S2BQpAyItFchgmm
A9gkj5wstuDQ+mJQ3JKH3VtOZnsLUmODiXPCCaMiXqjF1nUbjTLziUaUGX76SuUwIbyo6NOgt5sg
JXDMdpjIoEkJwHasO2ryZ1g9f3zklEG2/XpLc6mjSjfDks7zUT67czsBUK4GKOrikLg3pOz3DlWE
MJod577f00Sb5r4N1/TNNkrAauDpgYPj6h1GoQTbE59mc2Hswitn0DUabiK3AUCS1R8QMXBvZDCr
xDsBeosRkB7MooV3kA6qTLkqM7bWq0YU8zoISlSh07XZLYk+k7wADmZ2xDn5FCLmKIoU7FzVn4zS
JVb95A4I/rNW2Zni/siw/dJFbpS6VsoQ4ORs4CPyksbdXSdmSMFKreXZUU/UNQsy3XWTs3WJWyJ0
/TgTVXGh6Qhgs7L50PTHG6vozEVgrKO9wKFk8wCSGOpzWIvYW++rpF2FGHZaYLit9dRLpa1frzkW
A2mH26LNT/whYyLtGm7IeBcgCKz7OODmCYsCOxOiypFpZjnwVSbpb/RY4Y9CxOFz0kVLFr4JANH7
uQ1lgaleDt+atOqsWmnPJDUDXhCT7N1kYquqahq+dXbAc4Zywo+jjJqFydE+6IxjaMTs2K2q5mQY
0q9RduaOmZ6YMIFd3g8IWtZ16gZgYjFPtQIg0wtv2VjjXkftYoz3ggaErdDnELTHw+Rdwdg/1Gf3
2XXSvpexDQhdiN4CkwC+/NuDO9UdCfTwADuUx4oygOz30fnUqu7wbgrlmjSQklXsq5ljy6QYHjyr
LZKvq5evuJsey1Mi0swrcErDhJrO/WJSvL6BJQtkVrHkjIQ3dMQBFusK61AvoUCvaZSY2FyFdcWO
df1hj6ERA+QBiTrIlyISifb3s8evd4gOn6A6PrLENLTIyX8v3KRfLE8jshYQsbrsb0sqx7tE+6Im
0nYtf/vZd8KB1s0wn7rVkrPKjyZWs/HOgXMIDP84nkdWSoud+Nq6jRkODq4UinKBzhF/CXMSQL3f
yKnlf5WH0R90/0KGuhLvUG8dvyWAAO0M15aQVCCw+qW8DbYwzg7eqqyMXxw24ieTT0uS/d3eB/fZ
b0HVLwaQtjv7tUw6kzgtL5WBe3xXuyvynMYnPoY7Zhg0xnXtVf8mqWk47Dg5qFsqS/kHji1oRByw
v3N9Q9gJiJR/UYv94mdAdRb30MrUkDhqjLEXTonKZxTlIjamSdtEfWhdRc+LPwnLCWlbz6Y+/qzH
MvyBHZmxpdpFCHxkWWVKpAOvSqtkyLN+hiLNh7k3mHFC3EHcS3qo+tzY35GKLq0MItR80KzEy9dg
kUxHH6xhfciXCzeaQqmTw1BYdD1WJcNth9uoWJfyz6SR/W4HSJu6YO32S6L9YRjtea5F44oKSyDF
BX9dblJV/xImsz7WZ2XVxdf7brEX2Pm4b2H+B/+tjXVhUqCzH69DM6z9Kk6LV2eFeJ3Zq/0fHUoG
15xzxfAOobWehJCECGHGHrnXFsP6oiuUl7rW4rRVxlmH4NHBOs2ZQsMs4ts+dWNuAQoCINaWrCfR
JfSVem2AJAYz5SAeLfHUjLsZco0qDa51rxWg4Oo8lRjneVNaXSXvOlD1ZdtqbrJbc5ywx7Bx5d68
nWhORpgbBMPRAa+Mcx5h9bZLXpZNyrEd3s6wxXRvZD1RE+Z/d4+RBxhpXDgxJTF6JZ1aNvk1B7vb
dj2CzDNsKW7rpg81LXq9aTopuN77yKLKFobOG2OQz5/xhBQMsWKV/5jpkVbvrOmRTSVMY80LAfXm
wdOyZPfRDZ9PF8yMUGsd9OsXx6mpS2pLiL9uloQeifJeI4sUOJTfZcNvmbk4z9TBqBvsP8KWY1Xj
QjwxnBnBKQFe+JzckjttmMOUUkLW30HP8wY+wuH4CUI6wxvIJ4QXYtPEy87A6jYU31du4RriYIwx
3tsLax6IXJNlN6CXmyCsT2t5cyE4Kp6BcqThqn2Sy1fKyJBPk9c3HKTat9yVOWr5qLxZCd6pRAjH
bF5M634SjfXPE/3zluoGBjwURe3E3vjI//xs0kOtGx/LWy9jSY4ZSSifUhV1KnEI9MtIuKMYiApJ
c6qsq0ZPFvrWoQthsvzfKtimOF+J2qVDM85nZTMEdrPwi/sk1kbu/QFwEMQm77x4O85LKcLf4A/I
k87BG+exsLugrfFTpJfsytQum0k/ad97NqTIcYGk1Pawj3O0smxiP9OJCrUYdnycTlcN3UnvqjC6
bJq83HlWKZNOrHK7vWe0n6kniZqYrSpA9h3mlVyRcFWYipAS0WWKd9hkX5RzjixhyNjIXWtlpER1
Uv3C+hRF6+Ovwrjt4oH5MvmgeFcF+BD/PF5GsfsqVvFToVxifbLiQ7dsXgWoO4UI5DuWOfmfjPQr
n2AyOE0J3wgwFdf8weAkfkLbAeh2pmVy1ZH6w3yyC2iWizPFpWepTo+OuNIvM0UvEJBYtZea0AsB
mqQB5uakwLz6j9vLmzyw7wog/333d8VPrwya2GSlfxzaLzOrAzR/uISja+iUgssWTkgcNwWcQ7Rv
rzDycGoCWAPS9RKK746OOjOUclEXp61hiu0lhMzBwxHTTTdPUUVqNaNtBco3Om9shmiMr6wtBV/w
84jrnCf3NgvAQ8Z8qi/N0PI6uF8NPnOVfm9rVVbQndLKtKGZUtx0gpwe+YAtupDHN2JsnXpSjQoX
Pih80wEL4YzI9FR2FmgAoKl0Hcm3/ljColAeGZeF/UrCvXJfDP8lgx2lcpCFL6ntChH0psHBwhyW
3MIZ0GS/z6MHZsK18GLywJTp63lhdUqHBphACfYU/utfl8neI5aK8TElexDsA5C7979xyS0j43k5
NfGhWOkjuWlTnNqUZPvt3x1DXaSFTfulLqh2h+u8Sw/JThw9SKv0QFwQxsgS0mqv8Dgj1CfCOyEQ
2r8JK97pbFULxqJ+g13h/4VqoAhdguLHfv4k1j0lrnWmti/DrmcdG6fNbCJwPTF/B5XHaWKfoFsP
5y4OtET4vYU6ZxHIzz177s7UCqluGBomh+oQglYh3xG8UXbZGNf32mE/iVZRBlXk8lTOe3jmqdeD
U3Kxh49JJdhUXTbwrrXUddZ2X3ifKjvj6uhwwVq0ZLP0uQx42x6a+0Dq5tRxz79A+WCVoxG3zTwd
hMZCfd4BXTjIYyTeHewzQjNdxF0UaWPW5gsFIORoI2+FY8QGHrb9iVOiJw1MJqbaydtxXfrnadvZ
Rn0T8OP1qymIe9G5W9VTGRyD5MWIjG4gx6DQxQPD8h6rlFX9/4SGcHMfGo+lucd47NpVDM7ZdU22
5HdhKiHXZvOs1VG84OQp+NpbSGH/tJTLXn15vPVpQebnPBBqk1XUOhq3q6rcyLsnuzdfut1zDG5x
f1Xp0DVFb55CREhYtxT0FpJfBiokP4WUOTp8zrLrAOHa72pUEfbtw/tCAN0VM/EJ2XTPc1q9dH8x
uo1gN3mabyjnEehC71GS6C81KLLOLiLehnGV3/BXl3BkE9WsxL9dgZByE1RqFdpHb8LNqk+fNfCU
6pYs4LAx+46EeisOwHaf+YW/QGCeHV5NGpmUqFYdOMYo5PVpne6FIU7CGHvB8Jj5voXGaFDMBl04
ozKgfnb3bfYusN+Enz+UNMR4VzLJ4c1Mv+UBHA6sLAg9LGLO9NbimSmw8MvF1r2BL9wgDKlLM1TW
I7uvabEeLbe6COUkwmi8LmZ2WRgu6n6a1m79zxLXe0jJ5UJBS9pXgL99t/rFRsE2zgPPxDXe2sBp
8X1p1IoDEL4zCPOp4w2yJvVgz5VMvhc39lr1AAVoJ/FjkWkHTt6zzQNyWPB4YEa/UPSi0dwd12CE
chD3iQJCMzfXswX8eb2M7GDnwjLmWbOl4FAnpRxlbG7p4tRBAA3RAAtNDxDILduqAPPJ71ZEQY4k
mYs8S0r6SPkg9g7ir3HGdN8wSHOeNEhJDcTa1S+LdqcAOw37+kgfDsmGsYJ1/T/h3A10McNfbbV+
uTUeRQN7DACIBxDlpceKWHxTf8xFh70XCql0I7a5rUoZLZNPSydBwQwNYm0qnUrJoJnkxT6/O/Aj
EA1rPS8icRtxOXooCEuh0o2JMpMAzMxK2gL5OcFAJt+4FWoT4Bo8kpiKCUTzP6N9SNjNyDPIenKr
k0wYqNopnIEJk5L1rvD9NfC5nfg24IHxaCfabbe5aXZFqb6F6aBXUuO042oUqpW5Nuo3HB5IFtXs
wjut4s6chw9hk5+tRTVbOOCqVWMRk+AoqeILJeyDVYcsDLvHSKXjE/oitkIgeDqY7jra4guvcGaS
FGU4QAVuE2oAe1oJ4OQp4522sMhOzF//m4EdxAKLhJiMin3P/Pt6DBqfp85+AH3eKYJvAtwnKDTI
dVFGMApKEAbQfup6zCcx7C+2lRxa1LoUJsZGlUUz48WZHSv+1a+c4H5u1Go3zRB1WbekaPves1v9
Kq5jRFNoFvkHA8tI6cX5Hsp1vKkReuROrXSEJEkAXu3s7qDdDRT7PLw/p8HSW7bpBGo5K1PvFgUx
SX76rUcQQsyIFwsx6T7VSE5JLD/czQndQhS7Xhx0QYwrU7JGjQaWwWhK2hcHK++abjrMLRySKXtd
RlWi4K0jvX9oa7QWQeA6hH2KSucqaKssBrjZMWV7yLQGIjOAZZMrCjl7Sqj769C9T6QG2U7kaPzR
/IpiDQ2Xx/oQcH4M+H+tkcd6cSgLPpuJ4rEKvEIJmvAJSR+KIqqXT0Fi5kM1ArG0rEwhQxMnQo0t
pfrWg3Des0e5fr8qZpcQlmG5CvroQ+rjnUvfy4SqkiyLf0ETKy3Qt15/P3AJ6MimP97bdQrcQyun
b2nYhiNbelWRIVYZWcTEjVIrcvXCONSRD51e3d5tqExnVlUEyonVykDqUVHlekqeRdKNGWCfV2IJ
HTkwo3cAbmpiaFyPikU7jniw0TKKGBZaYxofG8ZbNyYoSD+A9awOLVUn92LJ4vTwBiWDOk0806VP
/al6kqzm3g9KZXcmAq+v08z7UlBI0fRCMRJ1C7r60659DV8P1JjYeLwcbZ9yZMfSUyHNyTm29GEH
DG4P2QsP72NuRR9KF5JSaHTa7OfDD1GiVc5RqfzZTu91+W4q2Mm4CYrhHSjj7hjAfmtVioBrHWYK
9alNuE9enA0D2yoeCGWLn5Jyqy7JyckTA2W6HPEe68IWFT84wgvBpT7lZkG9Spz0tgt7uaWViR9v
kVm/hNo7ontg0NbSNkeAdGlgO1NaBgBrCbzqc1o74MTmfh0YCWBdOtAWTy5HFddt0SKXiQHqWDHb
lcQ0Phog4biShPDh9HgQ4PcUtkVa8oZWh3GY5gFI16bjzd5AzeM+npQgTityu5LO+aOT9pbxAi9m
LZf9mlZQYpgIfflZmUofdqiVJjAW60f74xxNfAI3xt3UuhGpxNMHqrjQq/Rifh9v8dDlGRIf83Qk
uNQ12JCHShAultsMTpNS9vl6Kmbd1OuEhhhFF5qJo0Mq2YqPeZmiFhpowNPOctRAZTWg9LcANaJ/
FFvG5E9a+t7q16Jgqq6Y1dRB0cza2FVeB9nWnQV8IK+l8u7W1MXs7d4mHYjsWDFjPkgxAI15ybPA
uW2mSLtSAHRgx3KgIIX4dfIg/95JDrv1bNgk8e38orcpt//AZ05hKbABKcMQe1y3XTnPMyg3DIVw
3YsVDSxJyohj6L1Vs1E+9b9nuRSXB3OJDPGRTmQGRzaBaOpwXUEEQ97BmTM/lEftOTR8QkZehhyO
jIRW8nozgKg0EcDPuYDcFKlCmGi/gZw3Mp/XDuwbhfElO1gjnk0ful1ZdJ46P/X29FIRwXf9sgXy
YwH61a1+0v0yh/HbAvfdAILMwkJmtpT+4a4F+WNWBPkuvscO1AMwB9f4/WnmsBsHUr5wEDD0wPzp
YEOPJ1o+1IQ5Z4OdrFJ8yI4G9IJb91cMkw61BDvK/i2rLCsIiKM6GsCG1o4PRbXkiZ6trXYyj88g
diON3jBPdQIh4Rannd3TY4/nPKBwIyrwUDXHXyx2KOOCpI2dTB28c9v/LuG07YEC/MqR2fgit6XQ
ZduFU1cyzIEAqXzGlL+LbejOY+iMIB4ev/8RXE8Pz+oe17MghCUf4eQ0KT5tbJJYGVN5E1tAzDVY
bOyLUEiyWyU40PVkjGz+0VV0ty1oRpnP6492FLBWBXCz6JAVdIvAwPez8yucoxY++GXC+v/4kIjN
0kz2BBW4Ecsn7kX1VCC03OZ6wctrMu+3X85PgeWCfa92viFO06C1G4nxB8wKd1gR1Fhu06iImJ4s
Am0IJ7oDKuf2xBWvvr5gd7yi8w3ZXC79v1lUqwo1BWw04A9IgxDUhzFjHsdU69lxqRNW8jhZ+dJ5
PRfdW+eq1H0MW3d9unZdK4EmUh8Fd3R2XDYzFHoz6koW9fe3GM/e3BXnYS+F6JvhUE3+ms6Lfkt7
4R7AhJvdarV/jo/PJ40nWdvLnxbw6qABZeMarWhXRDdiwPDZ0Gc5UHgNGVgEOc2z+sOrLWQVfuYW
kjbhxWfubVXUExqv9CostA19MnXRrm7JCDZs73IqDDVTMHtpUsIT2HHBvXAkuT3mWZ3VoFPwxY1s
wcSrs26t42OgAXmG6uC2Uvma2cm/vpPLPDfp+0YjkfA1t1jEWhpI6exF3GFC5E92El7lGBCnQ1LO
aeNnYXvVssOJJo95TSulV0z6bPLhvwcHB8umCqrYFux0hnwQhBvYpOeAQqGhOqpLu+zGUWUxkEBZ
TeDceDKbVu+O3sJorprA1Nc6Pi+Ap/5gLHkz+ehDrYBCpUIw8hJ3JIWZHZlsf4zdpSamPADeCScH
JpcgrJm943MRNZwPZfzix8cwyE4vr9UrJHeQyIM5HIywKYsLTiBo6sb7WsVa5fFRZ5PJHe4/dqFJ
a5H37+ckrn2moTXKzBI8rZOy1S+K6QieFiCBD+e/OfeJYm7tLQzKKFl+iGt7pOWqqJT6aB1q7kdo
31wlBJhDRFfdSdRzUMj5Vu3wjr8p2VpRFgWwjY+rY5BcfZ0XGyhELwIvDW0aXKT6lKIxpIL8mbs8
ounYgTxxgIn0rHrC0SFz8YGxaqNSJ38K0S0N0v4x0lv6my6TABaCgJA6nGRqjJhyilQu5dEHTydG
0Lgh3WsGdPD2JoJS5tRai94ntNSSbMIokhBY6/TGbxPgkzA7EBlnSRJ8iKqx9HM02B03s23igY1+
ytri64ezMG90P0cY3eH10IjeRVievtz43HtD/EApp3MXsuRxx94zuQVOuKG+o/uoDqDvqtG0eL8W
cqUC5eio7+LjuSliumQpp7NigfHQ005+0FcADwsr5s0aoFlsfvyL02POTm2Mv4F7AfuNgiePxrSO
LECNnC0XeBrcuquIHwYIopyFD8bAn53+yPCgsQXu7gYO26lbu35F/X6V6lp5bzDSLM5sHB+rh+Ec
65BAc0divsTQ1qyEcRW1Cztnq6donsUsIFLpTC6Aji1bj0rLxInL4FQIIVMFk2pgegtDqCHrmEUv
Ovi4l59G3jZxVktL6XQttSz9540Tkx0oyfQX+/txj6/D1K3N0et/SKL98uc2tA0Rgef1dHTDUSm/
w45BvddMlFNQN1kUtZuqAsZFGiulV7uxVHYApb3VHtXLebk/MatiHDWp9DmxkbicOPLRcK22nSb3
pHLdYl02JrEcgtOfi/x85UNbzNJOYj9/Vvj1Ax0aYERdcTpG0u7OuBRPi2fVl/hVqfI17ePTzZxt
Flo4VHZ/GmOjCaSQ7zJT26Eqf7bqWclw4pz9NnZnHkZKTS96mfh2e2hT3NkNhS9P6V75PYesjcTn
Hn8C4ve68n6VszDHJAoE2vUOOEG7xo9IOJYiHDO86TOgwetcg3SQVK5IBWIQWLROUXWXNnSSJm9C
w+2n5iHMk+LWU/ykoHZbTCOIrl+dtLR1A2fm6i6uSpM/7YBcJaDE9HCxDGkYFsSY/vM4hHxRH6XI
rbBBwTCXRbqkJZMprCSYXS7FGrFLDDy8WH3PePZZlPaBFDwCEFZhvEh9dsE75nb19KwzRlY0wydZ
/PopdSFrq2ZNE9NpeA1HTG+OSMO7xDTRf/zLTrEPey0LWU/d1NDrJdhbL7WDExTH216HnGniyMk2
aC5iuJR07rhwCWf8Qw5p1gy2Cj+1s51YjtENowMsDzasPwDJ2LVm0NJ0s9rVzIuIYSMp7ewThAOE
O0CHNJYOIReLF2v4bLOTd2lkguAzjBvV9BSUet7oTjJo9OVucX/eB9ItH/SAh9c4EUf5Fv3Pdydb
tuT+krU3qAvnpGubhz3F/apfnXq1CCeA10BGPvd8/qRdph7lGnSIoW0aAVpf7kSsmUCWUEphp02i
xRXnChzzqFt7Gwt6iB+a6ia+Rm5zWYtbgLMHAMOYJsn8uB3cqGjDp2uzEmW3wrXl0QvlTiyZ9VVv
LCS8Rktz3ueSWr5dlh3UEuZY/jUmY1OSKW6DU4wMq+bokTgnXPEQjefb1MvSqE+wqcdzSoVoGStV
QNEFDhK2ivEbBdLGt++9zwPcnyQa2u1KBGChAAKREJOBJF7i0xvD+XmabpEX/tQzZvKnuJTwLGnm
2C9qVlf0sauZz0AKG17xkq9xHLRe+02RJZDaLtro209j+1Uu3Zd7mQTctCuNw9xp+E/Jr1v7bFQG
OB0Nr7kao7+4/nfNHOawdDWXhNctHoRCH8gFD/7TN1XS9nexpx/TkU+jkfYKSVjxZ/LBco8uhn1n
ZgZ2VJIzgb1F3Q8DM7TV2QqNQzELbkg41JhZDGCfOIXyEXFQ/Pe7aiXcWbUZNK3I862/evo01CFl
M9rzGjhQUvxpHceUoF/3tfxAH/qtq3D+qi4vmQkWLxVcJf0Z3WPm4Zd1QOXFEUfMgUGyxs/CzJx6
1DSKUR6YElt4K9ZMiPCkP/rmWkCgeiYcHQ0vZX50swRkNL3H+5FaR8TE/6BbirL8vYeBA+mqG6dc
1qz5UCakLydgaiIjmKK3Mu6UHKqS0HkCqbdP/SC1KxdwZgGSCKPba2STgrnNuhLAC9JfxJ4ZrjYT
nrgdELfHUIDYjNhGkXsWk/zr8UCONA5nMOu8LhIO7YO9l4ouhZ421/qi9gvWaOi1cZxwJiVAK6Ec
ADKD47eNBvUxhxeRiZHarfjk/K8lfCDiJZedM/EGnJrLSdeexUB/jfowBJOIpcWaylP120oe20OZ
V9TpgyeZWM+VgON6oqHfYYo7nfPJFXg32ytL4ceJg+M18+ETVlii+/E59gZZrr6MmxhKSu6JCO3l
+KN18AkYjsjMUloIdvkYGmboRrBhQPXdQOjnIBsLohdoQw6utMLPWPLCt9oTnXSL4p/6EAxaSio+
9z7M7OPPX25xZ/kDrc8J3W3vRPLja/VEjhEqETLrRx8TJAJMnISG4CdnCyMnVhrh69VpUT46cjoD
3fMsZ/4NE7KFQZQsFT9X5iV2nUGssR0Wh7rDpSFqOChNzKxgsW6JgNoY6Y7YYKF+tXG5Bl0tp71P
3hKunU1rkcSCdSrCDhAVXaZNhgA+dj/eev9OV4ZAfE9XjrnFbPWGV9w3oyxGVteML/scmYGAHmvF
i4w0s+DUpKXNcBKpvmLQS4sxydlp0t9ja92Ojuu3WGpa7/x/diuUn9AMOCKY/8cgNYgtVSAfoAtn
R9w+zGre6Fstm1WstjD3ywHM6ugcM/06lLee7iw3ftxglmoDhvt1OCeKmUuOuO+72xkHgSHNqicw
8dBDxGTITlMAQ37J8OH4U6eKWkWRXalgATeDP5dti0Lq8VnoV+A5SHf/F5QyM0sAKEtyvvVPt3/M
Wx2g7XaQs2qEnmFgUltQlIrw7nsiVCFFA42HH6s9uw5cWzEvLN153SEM9xSlesbB93jkGWHB5ser
2g9J3wPf33x+YQECC9xN+qA0CCfFU/UCaL9WiDBMSDQj/Y7ts5nLEV1E9tMNpiGIHNoKha3foJ9F
QukqJzap2rWznupTjSPl1Va6Il+DafbN57VT2MZRc1aUiGSzjT9YCFr5RJgPOUilG2kp/sCTF7FL
dBx7EsdocpZKzlbWqs6ug/tw9P1Xbz2LoKZs/MyFz1Kv/lpSgLUoJ7WU2kchF/GaB6jbGOH29ZH2
LMdhAOffxnUt+Hy3hjE1i32hWfNIoh3vB/RJziITP+Q/OpzZo0jltzqcDbn5csoxjp68jJRR2zSU
GZOjXqKsG1YBCXDUAw/rs/8faWhY0S5HWp7G2oteRMu8qf9unfo9/ahIZa8S2GvzKjRj/gWHVVJz
28dIbHtM0qIvgIGHh16fCvXRDl/E9Cf6zJEcPdlrJKen/slrL3XJ79lDp7Kkac/GKv2Dt0N0Su7c
ah71J5SA595Zp7jpj3UeHqdERoLPmWOzaQmkZWiuMBIPAxIOrW2oam77aMGjU+2HUB1iSp4+pT8A
aB/K0xkWpYb4ViuVgEW4VOQn/ZU+8mKIy0CdeWriimrPanpCWB8OMo/QhY8XtXiyidr7g1QvWDZc
aJIZ13QtJZ1OpKfM/ztZeQ2XRB8rAIbPElo/NYmbdd8nxuGoy+/8sKTHDgXTDcaQWG8Lw4E2NxZ8
fbj3dLiLnNYH1h1+s9j6PD/QRLKZbnYCWzPKOg1MxuUdwCthQxfvfQ/EoIItsaItRN2rT11Bbnmy
W6OOVKwLJSUYH6dEUzFM/qUA78kwLk0XnHp7hakS0BOedDirVpXDgRjAmOrolGRvWNEEEWxBSiEq
lhtP/OvGHTs96tWJk1Sm3ajEYJ51DV0S1VRYwPydODWl5YZEl7ydruAniv3EGyR8dZR2Me8R6VTb
kb2ivJ4V3hIYH85IBPDVHxEVXf9sWeyJQtK8ECDKEmJizCzifb8jsN6VTNptqTeWhLHT8govZZ91
XtqVg/4UpVBRQF810lrpZKXlPXrXlZ4qbeFYxMUpbRlwm+m9xtpXytdLfmJuDYxnP4JFtnIBA6Ft
24Ew616VjKXAawrl31GFVt+Fk1UdFanvE+KEGxi/PnrrfXMmAQ4tTJvpVaQRhITYXKf5tdqKPVEb
jiPiMlEWLPIUhd4jVCmjQ4mXkfpQnEBmcy+kSoxUw3fxrxJpTKUYasWH4O9ADATU4G1pmFe+XJF/
zKj21Et7FLb2ADwm0Aew2gRQ6HzDIfw2E4D1hupadXI30s7YBveCdL6BRqso2YpZrsutIUPAWifj
Mlvg7+nfTWy+rYUhBvSp67HikZ71zhq34EOxLwJr5bq87Mb3W/QiAKiWwKYpSMR84nFl6eSmLHwF
dY4MghhfUKLpd1GnfQ+unKPdphTjB7zBCG9KgLNdkynIcuMowhUQwbYeF9Q90AdgeXKjfsy+HtuC
9o0eCBjfXfEZZz9UmkHIboSUyCNDgR3G3tRg3Wt6lo0ayYaszBPfQ632MrHo7pcQ7jbjuVCIorMJ
PkgdtrAUIo2Iw1hDkXOE0NGdYwuyhg/WgbQY2WssDRHeXlWo7bAN5MC1W454tkecSVkCS8wvY2xX
LtxAuj7zbYqDla6w2lRFR3ZQJzdXHdU/GfKjaQh985Iv5b/qIRJJLYesf23A1QvDq78hwvGTQOMV
6HXH3v3gStZ2CcT3NssfrapWhA4wcx3KIjORic+J2ywcf9WPQSpeYIk9Vuy4BSeCRjcosDeEhT7y
AJ6i4tcOmZ3MeMgtQZFUZdgYrkm5rpwjfYD1xEvwc4in96zZwsqo+MPoJo1OYH0mK47oEe/I3mua
rMwIePnCW55wluUBNivN365ElpD4eBqID5UJvqGUCXabgeFQti2U3wI36zeMOZC4kWldZ5C0oP3S
8GpfQks+CIZ9Qb4cHA/W0a5uctLh0DAYoc/oHEPiS3NsvpVnbUUkjSpkwgIrAGV6w+e0X0a90amC
Y99ZaIt3y+TvhiTJtdsdslhejspRHF3BAkaTUd4UdW/+daC8b0VH9yA/ispdKhhS/cTiVSEbmlHn
tsjL+HwasK7FkDdwq/bu9RLkXRDIUnk8GVyE/IZohQnUzVAfx9p1gHttdezDzx9xgdfrrdud9DPK
vGVxHx2hea6JmA2iKpSl6+HVVtuB/n7x3ElzL6YG7b/yqRhj/W/NjXsj/wSbDu8Aqw7kULnil7eJ
blBZSIHqx0/2RQN9QkQs0MquGa032WCWgOGE9NzIJPIcgrb5DZwiXG15b4osJxFZ3hNZwPxVTuOI
TK7CZ7yZAGN/Ob91VylVU6mvtpylQX99fygcrXyVESiAnoi+0l5Pfrkq+rgFZ/81AsOc489sPOd4
ZVAr3nlM+CVNoZipfz3XWr7YS7MMkrfkGk1aresglzB++GGjCUX9LUf5TiG0ZVJDsyQzYil4sBwk
xjZNgMkMgUvfr3anZ0xGdq4GrjcTAHRtDpsnoDB0/SsTpq/pOeKI59iaGURlVQff39q6JnfgEXM8
9MO0dI7Q1Oyt9HjIOvh0E9gGcHMZlETyzHpLVAYcsBUC/b8ljCuMSt1W9hzbnzndJbgJHr1mvafq
Kckcq3EOV3EfJpNusrJe+Lg6Lyn8QTD+aqWAfuSTvM8eYJzQXdxhqRb4FjMRmrps8RaHslxLTPQB
Y2iACZ6nYm8pgwlHwVg5yw/pLp/da0jzGP2113D+sC9tD4V+Mc9JxQ0NP18NbaqThSZ16Bhj8zT/
7EufX9YAIG+7yoC4znGqQzyYviM6qDL9UcCmTquPYKGsoDbOXoYVXiJ0la+TfeshH8VaRJGoEWZP
34fCuOaNCcFKGv/n3mGfcXbun183KzDIIrr8U0gPd2Ktuh9WvuyEy1XNEhKgU4Adceh4YQKscygZ
m22S9kuPTUgvyZMFMCmB/iWg7uXJRjiMS6n7dfkHZhG0TGXollk2EGqiFEW3UwUz8v/TxziSIWgC
nNF+MEaCxHQcepRIDG5WfOpOIGFT3PwbUc/7HzqvGGWgxpmFctSIlMxU6CjGIX1XBAMn81KMTB3F
qXAcOQfuXpfV1LRE16zOsPh6m5YtCspwO5xwnUhq+2vKTt0EszYMwW8t6gQK3H/fBHTJ1IEzNpHA
GvvtaBLG6jSAYhNeM+EKU4onpF1WwUaVBIq47YoD8TArccS8+VzIgsP5cW1c6pIRMm4UO1ff9iK3
yr1zGWlHrhgZQ6G3ld8Y03aMSbNRrZGQjU9Xz8rSJA5nvM43TXFx5j1FMmHXOuugHYdqQ8MdAgfe
D71AlJ3+lPeyAVOlipsfZdyFCz8Vk6HUMqmgrv5mz35UZaH2bOlmK4xfF8mzOSVVZpKJqbR1bdAo
Orsv7wo4SqSLhdfMnfUw6mBLBa5L6BbSOwG2bcnvlir0ek9TsPK4VZ43uWUKZtzBvy4sh2tHgJo5
EvSEkITSUX6Ga/4gR19W8GHnVq58W7NqWMJ0jO0QF4bJXb+EoOKy6RqPTyK8t5WBXM4x5GXz6lgl
2Y4EZ/pdPGzIE6vABsMjEurfzSluM4ptBPafp/+PLimoi96lFJclr4USmld/XIpMFrR5YuTWHrkf
6XIpN2qNa7ki1Lwz/tfKXVybij0GXJAM+3Xbz5zOfKu65ofzDqnbs+SaIr+xuGu2xcl9UgRHnE1u
+Ig5c8hPLzWwgu0OWPKwusHowbS1pm9zN+6yTbAMOxoY6ZZbUdqgfu++Ac59kJzUCTjVeQ5Qy7VU
sK3NjZdxmXTyDepdso3B3IlZtx+bg1b7Oh6L4Mz4+xf4xIZvB1q3Q1x70m0dt8uJK3WaquTYFSE8
ouSYk7Qva7tqIF2Vu8jL9r68zfSUGxZf39DaNQSrKSW5brGHdnSxrFPR4FLP1jlNN3GzboFlanHs
cMwYicBc/c2kezJH3sr6H0GbFZRnJVkSHsszIw3NtaTrU6J7ojkjjVvA/e+fdwLY7gGKx0G5bx20
40rciI/AQUZFoqHmMpq1/O0yQXiVy8CmSJfM03HiJlaOwu4MaCP+wKerWcREGrI05CQqyFsax5bO
I8NWzo5rPIKwEjSjYV7yzcp9pbAFVbR+QRR4YEX+Kh6Y508Z5YxjsreNleYvexCsvcZ9D+vhkOEm
B6ubrCBA7jjHBqhv1AmuAFge+wbN7ygKDNiz5pL6W/l5EW9AsACaindRXWCj96DzeGkZEKh4n0Gx
k2EQ2CcZqKXh5Fz2mszoMuCgGruz7Y4+aIfaj9Qj+8yKJdprocSoJoVfqGqnUhdX5khzwQdkBA0H
FhZFGveosLZyIEgXJgLPzgOVS0RfMZsuUaA0FDBvi02zsnxSYyrnMUTItdBOp9ka2qje14wrKPQ8
dewttmH69pFLX/Y6wY5f1JKQJF2QUzu9c6ozf3KmoMqeNnPvracnuy45QsQ+tLpimr61VabGTr2M
8I72YLjwz6PP/Ju8kmyOf95FFjGa2Nh1ZW2KFBxofCMsSbONCqtILL5YDAIRzwx2ZoG28IrF4VG4
lEc5cek7Zfmg9Grbo5zGiWfnFlZpbEUeqrb8pAk/ECJ199X331FRha8c8AWcW+QndHeLrzYT1HQB
HnYZ8Cr8xvkciQnlGrqIoN4+zNWA/7lOGQ6PUwCFyE2MQdAl6BuXMdq8qGZYznQCleLdw4X0wifU
3TlBlTK5JbMbn/WLYHiHD2GpW7UMQlZ2/GGJaHPk6PkMM8pUb48QHhOmKq5y4tiv7DvjAoKSKlgr
NbemOAUMGSlb0G3gnzKdNykefFc97m4x+MXsZV/iFDLRc1YGsIzymGYhVji54Yi2vwwHMKZbUGjd
oFvZZBvRUyGqklY3+Wb7kRPbKdoMo+emqRsZVn5VArUhGmkBNTeAmjJLADgCaomQIIX7emeHXfVg
FI6aDgHtsYj6vdKiTw50ItpHmXm9bcb30YIGQ/u9IIClp0/vcbbntWWb/zYbw3QawAv2X/Qn8ipt
nLvq5Gssl1hMYKhc1DMc61bv5A2x3Ih7nkSKibTmMH3AbRenuuOXqyBdgFBR7GoN76J4SLPzUQO5
s/b2esNN1DeqtL2mmO9evkx71QJB/Zn5brE1mSdedGzYPp1SBMtPZp4Xv7Itdr0g7zFJZ4QTfpI/
KhmIeXeIeG3m6k/qZ79hWVBKY5RmcmFKJuFxuion+vqnVd2RbWfVObKvYA4jWkDh9PL8aXq5ahPZ
Nwh25RkftFMOAxFlmPrkSkMlDzAYhWyGKuOaYv1fKcdtGalTk7aSlSrcfWKQwIRqyn8igGvaRq2B
loVgbW+M3GMaPwBdz9gV7VqayUF2JCDiS3ofZxukKZJtw7QoKy7gtbmjIsfPbgXVzHoMDNQxXakk
AcBrX6iH8UMWqecN5NuuNwpxR9wVjkDmaAYnBA+tnmWjrZ44Azpi31nzFuKzk092KK8d+YOuuwrv
PkKi1G9Rx850oj05BJ6tqiohDCvOcXiLng3kPeXl/r28Hxa715ehKrOxLJt7YoV8R8Zsxe4Mwh61
hMNj2LZOwJofi1z0/HJRdIdmYLKdWkEAyedtfs4AoiuyL5djjLzUKmNijEjzs6AQa/HDaFur7kDn
WUA8oTmyhsGsX8XqzFbfwkr4pczQNS5K4V91Uoo7ca8vF9qZXHglzD08oChJr75QAQzye4/ruSTG
FgMO8iEIx0s0PIohc+y3DVUcyIIde+PJEDyWoawvE3/Q2d6TiWgESGSGdDPiDBvd9rbOHsuhnzFr
iG6HPTWhteq0vBoj4agwhD8eW55dy2llQ8YUMGgzhp95FBlW16DDlukMhBlkQoNi66gK8IplZrBg
UjwWDHPABEMjRuglNWtfypc51KypNt0loSlw2nqNxNgw5RdVHb60Tp39BLPOnHNl3n5Tmeb8D/fi
NVt4I922jALgtZqHjLiwxyXaYTVrp39NKDqMhEw3yJDrSRouqIvFuSvyfHVLFi0smgtTRo1Mf0OU
Dgt2T8kO8ytldu0Jg3HkwIDp4wBsrFkHmuCH/fDGRP8CwbY4whOKUzi2XmQRhbg6VHnyZwNu2SKt
i9rAHZR49x3ktuC6Bw0XYV80tFkFEF6phmIZpZb9hTq8xIlDZuKhs6cDH+OFcPJKi2s6+aKC1uzT
ZOapSYZscnRPBCLnSL6P11M9lb8tn8c6aeuz59NBkMFcVELr/KZ09hWr/L1ncFRDCjWwF2fbpkm7
1hTOghKM+BX2sNz9Csnk8zmWPThS0pZrNqnplOkRUJGVWz1bh/4nioT8+EaEZ6LFbpJUvKyt4l+n
hpF5kGm+D1tb7h51yGslelOUbTi7XA2C4VRiOEpedEFmZg9jWr0r8OhS/ATw0+lWjKFA2RK76OGg
Cs3Dlj7GnD3b/Tfe4ujSg6ftnqzfBtfxL1zpw/m0RbMq5my80yUlKPiL7qPsi1QT4vrWVZF1RvgQ
jdla17dI+nUxF2srcjLACkXM1cgNtXCHzWaN52Oq+b0gzfTVES8NXml/oAl0M+88xO8oUyyDyInW
G7mgZX+b6MoU0ZlDx1cs4D2j/iREXJEyhJCWpANf5IXuoXmzKQZMPZ8QhZa7sVPOzaHQo3RR9NEL
Jul7KtgGLxPURQzsQYamBpm9CIYrJ9ct9/u+wNi5AgBB5/gmi1XTs0QfwkPQ2oEU4bpJf50aqYma
v1QChtKNFi2qTs8UPjn3vLEsmHoAFvpR3E3GEiGavO2QHfQFv77Yp3KxCixVxwSBiNypw4l63Yv+
63ufVlPv7FswOuimwmQXLuhjA4FP6bnEOQ/KgGEob4Ts2QOMfFZRyujb2jjMCuMrvFlNftmw7hf/
yqQdB1rksuOxjv/l3hJmctu58kenw6oxkbhYQ3F32vqtgpGCVeOa7cy5N6+1Gs+zB9EtR/nDIr8X
OR6zgZO3x/CVDb/488jmeDn71rYZNTPgY1Gxjyf7gyaHSxmyI+SB4oUuoPyJQmushl2vkWhMnqVy
KnhQudn07EC2DBh8qXqrSiSgWGOmwpQSDNoQYVUXvEZLYFLQNFDCtIa2HDlH4+uQCxHZZArWd5vy
Y2a12CEkJedRIZfOZ5qzSGgPhtq72hl9glgJGld+yLGGZHWHMANZhuUVXN21IcnPxWzcxcdI9sUl
P/uqsUYUx7lII+UNnqyZJs8JdrHCQfzoc0PfX7zNINZFVKO375xvk5JyVxSZZwP3q2DxrIYUdMxY
84m7ooLF+Q9X8ntXVDjxysFhEnASAVAFpfrzeZiKL038DUWNwGCUuaUu708+dC5gP+dr/TqIhgjt
6d0eEdQTV3KSWqSW5STKyr4lbvUU+7ens7VS6PbbZXNcw+jKBdR28JmAsX0U3wMBUASRcISq9uhB
vMHEwyEDWI76Es10sZv6VKb+WSnfp+M34zPbCTd/wJE90+dVCXB2BR1SBdkzkh6REYdSnw3hkAbG
a42s50DZgMCnAlds5b2ij9klSJP5DAyYjkUX99qnCeGlXKzEWK/DToU/b044d7uBdpPMYTx+Tehl
evw4b6UtSRsurPgzZ4EEVr6UtWKaHWH4adG9ylVxivBMgFMQ3bgFB2N5aNQpJGT174jXiTLgHVy/
djmZnPIHZtJ7cQ8ZTurgFtZrbeg5rnfeWQd3fZk/HYoLqDngPrUEBog01p4M6JekOgnmUjHl87Bs
ZV2pc3ZNjDPyYYeLqJKA3qd5BSDbQAVC2Cgfa3dzIUpIWzs6VdwoyT1efQ/z0vo9hYJAhBIQBOO4
MzZrJSch8v0nRD57WHYTcAB/6dG6L78iJowu522c9k4//hfivlXB4Xg+1yLKhDdxmFDKZRO76WhS
UNWhw5gGNlMg08K9ZOUYt8rmhSABoP72sWy+Gj1NOOnLORdkqxjI5eIYTHbvxrTsnS1GAefmPXNY
skRg4Xney4cNoCnLN6DGtsG4uJu1XFHeaDX+ta0IWOszJEwlaNtHA58563qbSbQvYIdTGag/Vzdp
2T9kAKh6MPkEv/vEqbiX3clLTVOWkXVClhkA7PmoXzw/KYE4LClNxXJVpDkoSAiVxiUcqmlvyCLZ
S9yU6Z9crOVnl6AidBDD5anKvH2H+b71c0f8aLFO/OhTD7MNkm3BEVGxHI75zg746dXhWXTQDscg
9f2gF8MBPN0vEDdAxpm5YWp1PqZcdVJS5QFJOtxUPHzqogQ8biwTAwFKI6vQgttZ4jBK0UiYgKO2
msCduzCoj8U8isHCtw3WnsR94oZoRb1M2oRprGSdOqj9XRtPFcJtptWOH+sdtvPcrdIlsrFV/deI
1ePCm9OWL4WjC0pQMePDHDvTHIvyYW5z0ar28fX6kCXKru1dAdpgLVPyziw5j3iScQTGkdgznwin
wmfwx83olm4j6OSs5q2iBtKdXY3UAz1JGoFiscAnUXBpXMTzXkln5C2xJGwtpIpDicl/2cbHeDLj
WQ+bLlnBqCOkBCVog+Ftl09ZLFKDMqLzgni5zlMGkSGb96aG5VRjio4bOdqJzcGV8Rd8KqqMg853
NE6xtccMKkq29AIDCFjfOdSpy2O4+geRWMuzofGO1rzFSUBZLSLmQFd5ekwxmkH5hqcPcbF+LBEV
i+rjXUT96BRCFL1MOymEJrsBGLoV/Qtl7C9ybbhmgbu3tM6o7YO+HTp+SR6xlpdUIgzfH5Jlz0vB
NzsV9dS1dIuZRZrclC1SUmxiwbfBr+eO7bcbdVX9cuxBHSnwBbR7AT00wNA4U5/V13ysgpTeDhh/
86yFtPGIXCRZI8ZIgGMKrKAEfWFAUxita6iOTigUpcKpNHTWSo0WJ8trwOVY0TSHG/zqPci5rRwA
VZJz6zgEOYl7yxk9nidt7GiERv4eYa3Fpng9pe3ZNwRiTJ3KJu6B/AVhmnzPwbUC5claCdTyLf0C
lRfiJ6s4t3m89vX/GarSq2f1rd/X0SmW9A2R++ypGq5egfwg3zSnfnO9Szuq9Phg0dZ2fqZEMDcf
nBWNMOrqrMLn8W+BSCL+FNXNp9bpT/lTXda+p3SXr8W9+N1kWllKg+oB1Ez6LC7yT1tZsTDi4pxm
0TA8AiaI7eIAds+0qLnuhq+f/zG3fvEf8hMyJopWnjEinfsYe2kAnjZlksRCZLrKPdikbuXQc5Jv
jvqVjIfkzPMWsS7Ts3H74//TXJbm2lHkXcdSleIkwUBTRPeGlmRaaZsbRQAmq55svS9hOXLZ2jb7
0ZpFLeRqLuMmqq4E8880ufxP3B8kegWu8L3BDXp70vdiWKxFqoMqkPEMnykNNOFMnQfLQf0zvK/7
7/lEmZeq7eMlgXY0bB6GXine19e9dzm3nrbB2vm3yfm/6We9J9vGV0NsDh0XErGbMbZOyifcNw/0
X2zM02JEfh9/M+UVsTN2SLAFENiN85HAz8CvS2FFUIpqrnvReZZ9+UkrLPP63YJ6I1WHK+QoeR8b
4V6n4ojOL0CoiLOThaMmWdoAWDnhNY7bDZXv6nwqSIxwawyeB95MCaVxGHJsEQUrPB88GeTEzNFM
ybkjwgkMPYUmE874xPsgaoTHDte6s53jUMRP+2BySovKH0Kgo6dl40JBcpfKadhqypzDPgvi71W/
sta/MPgD1mfxacm0abVqr93AjtpiISou+eUxMM5Gmpbm2s2O+Vd3daKUn04vyznqtema8X21+RWx
JMK0LV0nx6peRwmGCOUANRBSQp4ExFZpMZFgG8IocQ9kMFzQy9PjTrXC760eicBTG8EodwQYqokf
prEDO5YHgWu51W52fOQ0GpVMYgNxN3gIegT0KaSrlA9VJqD1YuLarOBJKpYjTcwXVIm606LbTd6/
9Uo521Fj0qWDnkxHXqnwJIihplQZyuDcOOJkWydvTwN6dcFN5jM6Y8YfM99lPMAmZ7C00s7rlv2Y
4zIPbeVj+qcDNq57RTF3yZtFN9RhPirbXCZZYU7cFA4lf2S8ygOk5Enrp0B57o/h6Dx9PGlLA0p/
CCiuHf7AmGqIl0I4sl/lAezC+MFCJBgttTFES2E1wtgnCGWydqIv9bDwanRTQyP0Rx2EkZFDo7tn
N/vaPtQeft5dloASvJVV4ZgM7w6mDpdMUgwPUfAJD2lPV1ngJf1e3DCIjfhOyKMKFGgFBMg5fXio
8D9/GQklk5nW3meRyIvNaZrUh8sj9K/Ga8mlHfN4r8X6Dvi41SP3YNi0Jano1eqkSyYkKKyM2HyA
6cAX9VZhRPHzFq06TAZKQymHEm96pTqscLkcTdMx+YtmuGbVrianNi2umNr04Qz3Kl00Tu5uG/1h
wEX2Wja+TBUKxo0vdc1X5rBzhjbz9RbAujcvjxHfSbJijvLqD9quCFG35CRWkz+oZM+jg3ogqU3C
BJ4dWNWZhGSbaVdg9MTzdxDj/8T8JXozm3PzMWXfA7//KziBU2H5gGWnjaezg/tNCyOgnjE+rRPo
MqszpoteRVb7nWnm2220HYBcjQT9PvZ4UeAT/WfZTK4yRYUpgU/B7aQTe42abLrnakJ6pXZpkmre
TUaLfi82RgUnPItkEwA/RYgLpjeP5BvQYD/tqdfn3k/ISnWt8lX1LEwswqdyctADm32JaxAfDrkh
tpv0odkAngkhndu7UtEZ2O14kzrM49gkZpnHmNu4zLM4WDdMceL6n7n4sKmi29EF+h3ceXNEHFuo
wyh52Q10mLeZtqaJ6FE1qY0pa8/Z4GPXvOI1wp2PODv5iYFTznabPciCCW9OX6OZKqptuLj8fsZE
7iGeqpIfkw6VrA1GJ9PUFf/wAGG1SNW19jqjan8MhP6rt/bb3cz8sqtu5gSxtkBLG5/zcAjk3th8
PnM6727ui2HP5tkav6ZOYK+vMacDuW/x2fjyedbdWWRa9Gv6enIADqfwIWo4o/dR9WT9jjdK4fO7
cAU5+Jmp0176jpXYG127dhApTaGqHm/6aO5+F9fNa/7u9k9AYEudXiku0kzDJVNQgoA1zSEtLx0d
60Od49SdniMF2JsaXM0RtKC6CPeXJ6yEVeMK9l+Hd07DlgBLjVdChAMDWD2AUA4Gzzbvt9lGuI52
Rn9rxSCbk+nFi7VmekA5a81DiLXM8e9bJNJBVkFav/MBYvI/fS8Oi1VTLw0SEVo4NJlu3gm2bRfr
QyGL6ri3bzPCYRQoLFUhdy6c3hlhNsJNaPCCml9JrPF3y6igEkN9U4ZNH7HYgdzDCcGXVqxJg9uZ
gSmEbD8Zpj004PcM1nmjLCGZlHeW9d6HsC/xzqEbkvt/XaTlXL5cm4oI2r/ZzArz7cjkGcpkK6Fh
CZFHPVme5hsiOGvirF8MJ5YI/Tju4s3eGbfLcC6pHgsuuEKsMYMlwrt6fzjx0wchHh/1xPfJM4hM
oD4DH+l+my+vZeYbZz10kCZ+6v2bV0t9ZHaxWfjUf62C9nwuu9V6YEKUcg3hsicXKCfLU484oJMe
bd/ion5TngNKWnr/GEHuj5IkGyUULu0290zOeuMHQ3dxKfasu8z9BaAEuUctzx96XKDlWfDYsAym
4S2QyUemABVjRtoWOnObGFB7pAuKB7eoRWoid0M4r2vFsDBEdQlyiDnYiqLVg56DDhOtjJGtos87
rVv7g6U3HcVcxl7WxwLrskGOqoFDQ0qzAhqFdfCyTcFesspR+4SOmvNC0jZ06PLgxTAy4d0otvGN
XHb2UIXKZDDcGDV/eclE7aO5b8W/pFou4yLQn07oPff2nRumaOj+JDGv1V6CgrSBCZrtBNQ9rPQk
InIAnNyVODFLa2REhvSpJUOvUzHmmtJwKhoBPJxZkjXcZsK8xJNrJvqnlGIvUPDU3DPp8GS2x83/
ehH5D4SCGjkDJaMB3utPNg/zTQwomjT3YOcLCkL1z5wCSvjs5f91r9ZQQftDU1jeaQ3nfwmWppRX
mi8Z1hb/KW0fOqJnbf6CLUdOdtr1lOqR+opepmylnw2TEg8nfgye8qHm25leoPbGeEDF2LCgreRa
qHBTkhwyCPysguK5/eImSNHmqyLBjkjWmClLdmph/ldcUeIslr3FHeSCN5zXHALdnzuu1MY0St13
fMvu9t2lD5Ppc57VLZ1O7uMYwaXonA490FytfTTg0sj+8Lmi0lQZ1Uxr8PjipZX86yZOPFaGd5eL
mcWQBErVDe6MQfltS/CP/yInpdCjIBnke3I4RmT+zpoD4VPDEZ1gyqmTUN8o/4GmXzQqfT82dgCa
4e9M96BBCSYGKsA4jWMJaejPL/OfXy0Et/djv4TYCKhWRq+Li4PoXBcJndpQz9zFCPgg8Y5mu8vM
KV9BZYirxneOksS8i/KfSQsmGDOP5/Jj8PHZ8a1hi3+DVbtVOuIDyAvDxkXq7597sw0y0gPd9GHf
kFOmR83WEaqhP5HMHlgQAy70URqiNFJ7tXRtfZliWiPh8fg9lESMV5Wk+eqLZy+nkpYErb83XG5B
JVFHVyw4gURbkAdZ3kqmv4oJPlhsa/l+W17fG3W6zJF68Z6HR4+4lQrySc9zZMbA1sKFPrKUJ2Yi
/73NT2/7mnRtPed76eqmivoJU+iTvxV3Oobvd6A5zCPFwjuGfHs9JPxp+qypuYzpKjOHlhMJ4Dwb
VrIVJ3xiZrd1DlHI5ggIsr8bPPIQDr6tSw3CNmfhS/qmv1wxz3+r7M5Que+GkWln2jyN16Rl638M
MCpKVWZx2ympHG6Oe2eZEkgUxU3JGzqTI0Po/vR9CWWxmtGYkQl9sZaAEhbxqRFcuvqd+zb1iCAR
ME8gTrKEBUTJUHbLGO8yhLKcTrTalkP6bvhFqe+bfSkEgtGl8nWHIHAGLdN3sREd+eFsqFdxsFoQ
FKAeVY/VpqVc92g7tWoGuWL5OVIHljUsV2HWmKgX55BCYFIaEP2eBxrrfR/wTEYY3a3iEKYpSLzw
eXFzgB+nCPmKzfJAmXlr8a4E2lCDpCHNh3/Fv8P6i3LMo1TWWrEZFNaih/57r2WdIFuLeTjszQCC
m4cPAkP91bm2/QIJMzInNGWYwJUnGc7RrmBMO6d1O2vr9Ok+j6bpHy3QqWT00r/7Q9l/9zYFjwuc
IioZhmY2aI8dmyDMSONpgncBZv+LiXKrKdpNiduF3y5adreNrUxJB+TKZeqTb6/7pxz2TEgwJPsh
V3whVFhI+haeoPmoKz1LB0tHhgCO9lWwkULuVYn4kwv6VkA+gUr1vR8bjAS5c6r0aXxpjIHInSsb
3O8UfOBxzbx5HoBgbBAWvQRqhDQsZXN4ekMq1jblbGa0xxlXA6+sQ31VRlL7K2dvqUhSyMEU2YdA
OE/15sR8WLtVJlspnPxYtDQPwo8fx5zb4DAsHd6JqSEYEPVqrhi7W2SKDocZLhYXPLMBvSq5h86z
3lC30YRDTJ4Ljp4tJS2ZgNRvrD942apGICtuvBC0f50enLPa3ORJvqAbaNtu8NkkVpB/sq32eTed
/mSygyW7AF4Mzmof2PC9kNoU364RbarlxQD3slLEJw2S9an+vLf72xLsKvermCceDLD7Wc5Ucxnq
lDd5mgxm14gRWzbDeDPOlAJf8IE73mR60kWyHn2XJTtlkh1PIuoPFIk8NsGon9wyy7HRl19Qexg4
yFybEZPXmLWZOqQZ+BjEw5CNaKvhlzH3rh28Ll/25R9invB7y3Btbz9l1STQormroCU5WoUVt7Qm
MsKYCoDipA4iYZDGz2KeLTv6VpJ0YzGxzCYopWYn/DMUHgwo9FKyy3xihf9SXe7VMKWb4XlCfLeR
BwjmxiNW+G4ZaSnF+KffsEiz/xA7E2omuHYSsNMwmvrUIvkjr0wl9QUk9+2p59khPiETIoIAnKJL
TWHW+ShmB/Uuna1Li5UwyW0P37rnN5Y300wEH8PQyT/XFo33Y5/C7DCy5wpl0C5GLST2f8E7tOLk
J2CSd6gczya777elwIwxxsSrL3pUmjpYMPIWOFQ8lhZIjN6SqKBALI7SVVxXpkJQQ11OMku59F+/
WJXOLRsnN2Y5X02yERPddt3II6iR2oGvQhhoMosIXWhJ2N167qOPfPDRoXqUTc1yFhwHXpkc9wGl
Td+B/T/W4WODRhL3zjPf6gU8deDJqQwk1TyN8/vWIL+CNEP4IYZLgh92QdKeSB+IymCC/faZMh52
QcMs1BtxM86oJbK6kYoyMH2g3vEDKmdcFYSFDU664R734s0WTGZJIyFK3Gn7q7Y/cZ3DFTsWh+4S
zb8WFog98jFyEthcOQtK3fb3RQKj/38t8AUCHMguqbq3zYyhiIxNwgLPlig8pjxwlNCt/agszzSx
ZeOiKFkUdRZQc5HlC0cmd86N7EgpxGJDaVhZK7Ag/R3VySxYn4+q84yZI8lFH8RgY8n7D40hMQie
CF5/pyJ0G44WhklXtaoL05QeLnS2Jhiltz8NvpZkaNEYON9CBrLY11kamijkNWSomWTZZPYVap4C
1WBXbpfgnjxP76jekMvOIp+rGr4z+i6QqMUrZ2QJY84Q7UiNPRU3y8uY0I93keFctOeyd2JXfA/H
FhX05lRMMcM07doT9Mb4+w++2wSYV7dXgjhzKaI+P3lpzrpqzlIS/FhMVaTtfieQW6acVenLpAZe
r0ZxVnZyBOh6yoek3JXNrBah4ViR+zZS2Jk3QXjQnhpncd6g0Ih2d+5Kfj8XH6YJVf+aJBdZbyMw
njkU+96TIirdYuCIejeCuKXOe3XvT0Vzsnp5usqSu35cTpZUQD2nqUEvgXW17MMXLYoRw7dUN+Ek
4i2iRn3xZ1dvS4r277iM4Jnm1imI4a0V+SV5O6cYyM2K9f3z58o49OG3I/47LEGtuUDsEqJavHHJ
imNtVqMfYZ75wxBgXH7uSvYylR0X/z9ysaCJwQHrcL/OhjwaENFXyb6k5Cg60ZSrheeUJijbvEgC
n8yYNxF+I1s8LrUCgl9GQyZVjpxmhufcDEdssKkY+PeeFrcjKoRA4oE3vTD3I9m5KbGwI8QnFOBS
2kO7phk2aJKA9mcVr+jMgSJ4S7ikMdLocm6TX5/a/ZlMsm+WyfwRrl3Ql4CqnuPCYbjNJafVYZF/
L3i+8rzoHCdeQyS/i7eFqLFNnG748HihmOi0P++OPEQ1fRiFBLlYHpW+zHuJD+A/Wk1Ynvxwj9NX
dYEsDdnh7qYaQF69uzKFUVx0spjoPZAjIwb9ouy8/KaWGsx8FtO3i6l4HfgjwsU3wl19tMwyd/6A
8BOJwIjAJG6C1nZA1j0RPWrBwD24Nsnspz1z9HfvEPWxjSFVn+mvQgIyldo1sy/zmDDAQ3GgqF1T
5L2V7pP8fxd2BDIENX+sncceNMuknif/s6pGR8RRDMT6j2dOK1pFzFdCgYhx3bxlMRniKwOVor96
HFu/6exHeFej4D7xYehTi+GEafowcPSrpXqWJgKQMGPhd2sEOgGyi/16dtMOMwuFRCObICYZboWi
ok/1bxaXGIp8y02bCphNgTCM7V0/xIHOMs/OhdWM1pM0++GqHn1Jx0bQ9FbDGzL4nZeUjooilH4k
q+QkCbcw9mVJuBo5CEaqYGSVH/4k8MkrOqLSyPYsaPhoRSNYSRVGvLsUJpmXs/EpkYDOOaYs2Kpf
hVrH7Q0QcYoIOlJqdwiwahEF984H35m0kRdfFNQXS1C+IzJkK1PsiN+ubxFFW3SqEQcgeRNFCstu
n7w9JoOe3rj+CbNqIZBunQ7N3js206ifiJJb5M/2KKYP+LKkBOpz4xPrY1+ISMcue6lwxLXDEd0i
qLL1r4U0A4YTKlhDzYOgzHVO/c2rOdMuiTKzTw2a4q4/UhOEXawn/GqX7LEGmUeGQlYhJVmIud0h
yzdC5sR2tUwCqrpFTMw2dyVzUgpV6RFhm2NeMGSdCkUKwRRhd5FQoiZ1ygCMVhMkFfHA8f//QQOH
zchBUpmMwtJcaUvXz7w8UX4n6/zpvBKK3aa6y8gpkhhSjhacNbaz+LQa62qSwNDHUGZ2LyuQWK1B
gJC0Am1IF0/alM54ThoZjdBoWP2OmBjEEP5gfNUWAVGU62RMz8gByYUi0tX2MWFGbJi6hgsVRDHy
j3V4XXE3k+osx62DZoWSEVcFf9QcEp78BF8qeGw8dLqjhpnd2PiXzuirLj42cm0M4w7GLVEhPka2
x+vVP7eES7p4bLieLDUeyCkdpE2ZnMiSZY7Qdvlx9LQLW2CCq9sYSBjig6VMQtJBiD3MnuQeWb48
he6rvHYj94oem7m+GZnx2+9y5rkjUhgq4TX7e4I41f5iYWwVuVpK9rj5ZMW1rGU82eYE7zIIGXtA
UzH4KNLtduFA2c5Z4iPELVQuaPo/75bpoaSCpJ5NpACWhN9DUKnJSFZzfVOwwPqbemhm0UJuc4gw
h6yMw66rCrgX3p66zMKtqWl0JlSMlqWCrZHA6nEXHG8e0Yrm4x40uPL1VblbjWNbtXCs4IffzJfG
/CevTtqglkIEDB57G88616nLXh1z7FJjxrCByQKQFEzVEz8A1mTCb+2GqM9yyo1/jEZlJZy2bD4L
BqsCuUK1lMJjr3N6GpY/9gVOe/rNxUd3yEv/f3lLhc0MafuHKJHDy0n1CmHJbuUt4PVhqH694C8n
7kkxvTelOS3mxaPa5S4Tw+GEED4lA2UQHl5xVcXMR9736iqOOAZah2azwWvhhCFjwsq0NNpRU4t6
DA+FfdGDnnGm6SsiuveBYFUypCYf6HYHytIbipbjbxoBynZZNg5p5F6OvoxPscZFfE0DHO18fAhI
nVzyFZDDLoYhGYaYkwFtdO5sWnJm+JqLHFGGM+AsMiaC2TVGxaegkwFdUUwNQeFX+RpfzuojJQ91
5SP0SkZxdRE0OKIFcNpF4bZCre8vD9QQ6snwKYDHLN8+wOugQuuRV5FMMCcyN1X2BUcwF5Nviz7v
7jxXb8nKmutUQ/kadVZN1OIV1B/gzm2fWCZFW9AENZgUKCBIBkOPmF3w6nJ0BxqAQHZfL5BPanP1
gl8JEIZfMR3atOJVE3RvdsIeiGk/RG2+tQe9ImPLGT2NE7x333KwcdFBPy0AudiEVuaJ/BWIVt67
hhTGuPgBVlHDWmgf5YyIsHLZcq3d0SHoYb0vKaWpknbv2eJT20IeSpO8/y7M/5CxqDK4rZoGqSbf
/vioz5mOCtrdzrhCjLVtpqfESfMj/E4LQW666Db9DXb5s7dtfrUavmv+9kbu9AgUl9/K+Yw4ERA9
HTCrsfyjZXDvM4a0BN01qQWErFHZU019hbpiDI7fx09mGVw7w+jRF+8+hsJUBp68FXaHQzjyBEPo
GoKyFSQxDHd6YFWATJgi0JAWjJw+7I5jzMDvhCmPwca222TD8X+EZLZ1rOX/GOBcJETiFhwsLgzV
Xl8WR5kowbs2kFA0Vybuy6F9UG6bTZRLjklxY8OGCpIMhiHde/uc2GAMknURwLoNbFEiX9P8R1Y8
iIS3Sh6QFBatlk7+pXoAGG3QRshQGxbEVIFrKE4WNucjc/En1KcJDE1mzB+lC0ILCOTsMKrCs4Ip
gxZzQVCjVPQeqHXFcEonHXwzsCYTuuR4XisdfkORP8XN3HdyvPAcxyYUS5DIYNh1ke9nEmPlim4f
zYIUb94XKt8xDFOc57gxxcpAW5JIMzav1ks062j/5DqiqVvSeJBIPvlwIwHm/4rsypr5Rnkn3tRw
CYvqD/rUWOD927YbBJKq1AY4b+lSEKj3f+ornZTUaprx0N3miO73EaZZz2BNQ8S5kETbcMqj1Mya
SSImqRBWbPTCdPQQ/gHQE4JwqygIi/FItmfes4Z73iimpsaGnD+/jqASkclcmxKBreBkfrybU7jI
u71M2qK2Z/TdyvaZ1+/uLiUzZxXbkufUCdyVpj8Jq+H/TTSa92022ZAnQO/N3UwhgJOoqJhQCEAJ
AzJNlwhpTgG0/21MS8PROdjerhf2Rj62lOQD+NZ2Wo5w1Ofcj1nd+Apl5PIFANA6C/KhAZO4BAe0
LfY561aVLgO9oN4a4+/khEbi9LRabAwCVAq09UE4+jWXdBPPiGvdiGsOlKaIqEeYZfwl2x35bRM5
G98QsV5V3MG3icpqnMBSTKgLIL3Ci/f/D2pFzJqJzbbuvCqoUY+V25iIGAXnXfByGkw6oeS+zsf3
mkTPvOj1AdVILu5rKTJq9YplF4Dz7BZyjXHlSGlye7SQ/lHcsOI2XuEENoWOcyMubgFca1WvuMcf
VPUr8/05kwcLJHItgQsQGUkssNKZc0zM5HSFW1uWRSs7qm7jtpJZMMT+Z1fW9BC+4miQLv6MowG5
EUcQItVP/prx3QggTVlOpODjxsyQoHxlwC44Vht2XvpEpfkDHwFZoEcs0f9Aj6uGOTiBRSIKAolw
KumLiEIOO7Rd2yY0X0fM46hYaD0AsB1nRcM5GevlKqiioqHqD+nY3XD7Cay3KPLVgPHlqBAeSd19
dqnAxnKKn8J+mNl3/XUBxM8Cs9KFRcPOu4+sroW5OTkYjEQRN2NCN0oBX3an1DQ61xkerKVZd6B0
cooZSEh8/rpKRF5c+hrDcEwzzOqqFJjMKftDIVU1A8Dop2nEBA4/fov1e88XBgA0BUYO5qsuqw2+
kv+RVECIErXrHKChz+vEIKa9QAFax6ShTjvSDURHYYoqVT0U7xWiKSkUS0AYqtTpRmJHWzuLxlwr
7ZFzR9AqcXJO2l9A3Z4Q8plfrRMiP/GEEyo3zhBeycIxMCbrGVuz/Cp9wOwhKg51CTPzFrdiYsB8
lUlDl1LwdUCenobxOH7UzqsWbi7Ag1HbmFU9DJDDOl0WfywhvZHcEgEn/onWf9vl9IIP4dJ4qFUA
Q98CyznBUujUlYsWnqlwLCtpot9+TvU2duHTUah/OFuSQUJoP9p50FLyTxM1B/KsD9rwx9aTQGPD
Govm35elHDSrk1NuVL+hFrBmqsW6EMSLZ7HRgyakxvbWkNZxw91WCbS7aPN4HfGbGkxCNnLS0AEB
Jx6twieQ97jA4N6bCOEoHODGrlY8oQ3uD0bF1pLPZYjD+0x6YLIozN5F3/W+9cOfdS97z04OSRzW
pyf6ibD70Zo+09Y/EI51g234qwYxht9F2/cX6QWtCjIBE5pHIzdhW4PYP9vwVlO+XwMjstW7z4nC
3c5jby1Qk+kHO63quVmqSQ+cGkOCNRKKEt8RetGIrgAzln0RgQlWSlqrhezEMVlga9BCAKhrcl40
tHBjUA+FFfzyZ5Xc+a8NydEvo1L6lERXecxr9d8vuVPH1IhtqMBKzfuKHJVAwch0WgKjGJ0N1nxo
0bL+X+jQxXCdhD6GbPkkfagEHaiRYfXrvamOfhAZ7g/aIO5mUBIICcxuF5Iijv9ZdekhXQOQNz0E
L0H77vU0KBE/Htu5/KokvlQ1tuvggpxesuEsipAf7kEk1jcgdNICkFsv92ouyRR1JdewuoyfQDJr
oZqb1zdRBFOvFmZQ1s2radS/H0CBaKKu/IABoCWqDNXSgktruXkVMl2R/1+/Va6Jbjh74IgIVf4O
ghW3BqMIZsXG4WcRy/VR80S5CM37GEQiwKY7L5d9zxnxMyXfS0xQcJrWEXYoeKQb+PwhFuEKXrMn
YErw/aHd0N7OWleywG1g4x6hQCVAOKkfC1R/vLqqw5A6+0zcQfY6h+dku5m75/EyZ53qZTrnJyyC
aIss8Ll9aBsperw9KYhCNP11pZ18cQK4LPOvTKjelZuxyKDhxJLbJ6JYi6DKOzqsd7Pj9foGqBpi
I8t1hh0pebtjZnys11UG951rJTdC2L7k5LY4H5q4Q/05xHZrUcgldTkg0k1XofKQaY+TRZdnNXpu
wL94Z9I/0tVc0HzyEJLBOZfuDtfaUl2dzHjyYTCRrG0QXK8IfZgZ5zf0ZE4FCEKJK+p1U3AaJBkv
h8hhBuJTsyh9UtwXpePyWKbPBcbwOK+2/lUqrFcAI3CCLdj37dQFls6Me9fDVrUWG+SO29zEThsE
hv361OKTFLArrGohuMlsAHwSynj9dRvsXyNm0+V8J1RJwHC+8RzClL/hY7MwDlsDPdSnmkNlUSDP
HMNeEgvmVKTVMyE/270QZ/rT83xI6/glfG1DMRbXb5fBvW71CUPEXRR4jvvnmKTi0QpyIli07jtc
GcNnoOyFeN0kW0MdLHxkxn+w9juvXM7SUUNPX288jrBB90hsTR7U2p35JO0kYopbvU89Ui7KJlj4
Js/4eAG1yQz9sQBrMUkqCcQOE92pDGNMQ1Ifi001FMwvuW9FDsALDob5R/RYboPBwo55JtWO2VG/
zDwupuTdl/Or5bDl/U+/McabVY/C6eTFMcUcsVdXSFhQjNJJVT5wzoGAOUVe7liQOVTIk9lURByK
v4Y9sAM7rlg0+CCSxM5KMqCsZ/Zz88MTFoAypqm6YtBBkpxGfE3iF0IBcrZ8VRY8zlaAjVXHRc47
C6isrPYuT3rzDiFT/D8ixNgyouMEaL/jrIP1TfmcDu7UJWOkyPgFWrJ2FI+mPHJqdFoUtCmLEOms
jyV4nhac5NAQuozkth3K5VAVopxvxDSE4PddDNYa2wT6SyCkgb9oE34WuCpaP/nI8l0iiTZpKmng
3ZchIVjh5AXuqfQOFs/wssxtIpb8QzkncH2bPFgeAbW2ootptMjhd5xO8JRUgZjZRZT69fsIBJJf
b25w2NXPY9xZYWjzJv3T4XEeb0ThN0BK6s8d7X3XM90yuXYpCE8DeHOW5evloiw9qW2R465da2sY
LSpNBnptA1c5qaOjAnIVTHe+grRYAcjkhXqW53nK80xWo6UJAeCrPMYsr9f66ZKAVNe9sMEQaX4p
RtYyVY3IuCfnaoOVGQuODc2HKtaIQfULfDXCubRuxVSZPtGBZAmrPvC4hK7m5pV1Tir7S4N72rC8
1R4Fq6hHOA7jJshFpndazsxhXKZdKlZCW1jomPQzWDqRqDbcKlFuKpbgqf6zXK/FCyDdiVSvJ2eU
L3It+fnQrhXU3ji4nnf9gdT57Px6h9ntF+eEhTyHB0M41W0cV3ojNhi4W7CkJ67DrXdqe6BqGgXL
25GBg1mIcsWq43PJRmnOFa4yC6OJwDUnDuPvBC2VYOVn6B2ITcq2tmFk3kL/9rR35+et8xG7mh+k
XD12RW3YY42ahF65NsK6kDGZwXHzYbXKu4psDBNlpznnxy6dVFYua7WSo99kY24S1Yipn3jrbKBu
T++XdsoUsD7pTXPSzqeGjuUZqYCYnIGYNxZNOvSRfwOYEXg4OEHmOOCBn98rpMDM0RQkoDsa+T2M
od79oi33X1l0rh9gQ+n4tGltM6UvtnlcvMiIBF2vl9g0KdGe47BofL0M/rvlkcWBtO3fibX/pBUv
xvV3iyA8Mm0WsJyN+Xp074V9xfVWmbOTgHJV9y8h9C6KVlU/4OYela/5/UoFEEr+u2SSfYpUyj3y
655L5OsxpDNN7y9ht90vdXA9Sym155iT9F0lOjrvFsWGhjgedvXQ3ExU9mUysoZwrsifTxBXSpY4
k5uRCZpeVYNqYSf9F5Kaz//zQ25oyUbdUC9OPLuN7FSlv1cKSea6bYgeEVQ0AaF7pFdoPRGNxbWO
6J0PtU8ON2AyEBqNkAqjXciJHufDtZmfGBmSWOyG7AaN3b/9PLCrHau648znvAN2SCEnB1QcnX5Y
d3kqpq8ctrNwoPyP0HplZlKT3F8leqv1YQLRN4H4zxeYTXGydRVr7zYQZvthMV96EonbyliR46kb
3tSmj/yFXQv/cquAanlEX/tvCksInNPie2Kwl65fZ954Bou95zFgK5DKB/fyXg/l6EC/n+GUNwsn
/rEWEzyFWq+TqCeF8OnN6141uQq66NNLrniiiQflTLG8JNZC9nXpta+7T5uevhTZCXOS/4EBDyL2
qEnbpC2/cWBNkFEGDUX8mpQIrS49ZdWOSC5FzTlZURhtMaueJK2Y3kYUWo+zTPzr+acW64VAikSD
rVXMkdpdSDz8iJtUD3nCV0E0utO4hSGcX3OsisxuuSVSYl3AbdzvgB3gKVy307pvkxxQSfRXXcg7
Vifmom688NcYERIC6NxILpMjozcODopBGWs2oKcdzwNNfDCTpaFtxuIdiA0WQXZugokNHiSMYV8R
3420H6Dw9/wyC8fE2TCP3MWPtbw0D4UHlRvNhLcE2tYGGmj+T5qeu4GAkxhEENcS7H2da65L+4N/
kSOfTEhT7geYblMpOwJveg/vovVLyBcR6Z9grOBakxC48yiW0cDLAXE5qTj0ME3NeQ3DCGhrHV7i
nvNte6n1fodmvNcxMGIxr59zxS8hALSPhcha5NsfEhTyF/mKIU1CNncWe6/fVlX/3x29gnXQ3fVZ
qGNixT7zY2s1z/gu71KYUTDo4TckknEjrqQN6hom2PCYuGVQghIMaSHMunJmX/dhBKqp6BNR61L0
wQeJhpUMooUNrJMR9SfTToOkcCH2eSGNT3PXxr1gMMoZvhiGyXRNS8in1XPdD93e66ZZNnl0bjuQ
3TLNZro4+y0GdEHs36245at+TPcV889ymfp+5Pwx0bfx7pjLxc2WzR497DOK4tkcZ/jD6x2YeLuB
/uqs35G6tb3ozcu2nXeHRGnbRcHfh/50U+FoGjlhttkb5LZHWtqwRSjemog9RwuL6YT0wwKsjiho
ozx9jhPQPLejall9JyB4yDoV5uOncs4Df3VowuAmC6zYZ/hzMmni28g5atcXF75+GfTzeSgeN3Id
NerLsOAmrUgaeqrjw5pvOrg6viAm1UHHR4aM6tr9brZ8BbJUfDtmgS6EgYSVymtoyoHVTFusSrqW
gnndsFnQ38LNeiPC8RkQuO0xaun5p111ADKnVr16aI0BRC/cYHdCUI9YUFHN3i0ZziivumagVXj7
EaHQWgl2ICKWjArNlrVBWQRzxBbidKT7yKhFbFfWCj92do2MhebTa5VSDM1d8YBLZllNm03Aprfh
IwXHAaydRWCbBST5z+TKmIQl6ck7OXrx1famWwP1BaXLV76W44KOSzW9WQ5ixoJhpDr6813CLe4s
hU/qOrKch3VBKFgJy3BZO9cUgQaIqPLUyZfnHHqtRZ1+THHWpjKyQvbEwsoltoTyMAPQ3oL7pYoy
DZfZ5UnbISs4PSOdQe+m62eo6oiymmBiV7YwHXgAD25+seSnlZUvYzmeYmL+oghUpu2WacpIOAPF
bUgVQan1yi6bMdrFR8LpLE8t98SQjZoEf1K6+N0CS8XuI6uVa3RnspYAPxFfPjACZ9XxYCN/QoFO
wccurBSouHjTOvY1FgyIlbjnRBDyk0GfvFpwYAHQ1XJZHRIQ3gOlwc8vGwIVHSEL+ES5cybxEEvM
j1R//J12dasEit5iSPIwwY2U5KCRRBCA/BWIIA5n/tYb7dG959uHLvcUKIeBbxEN0sbCRBNu7SbR
ouqWJsxjEByd5t28FJPYlebXk68rPk+5Jbd53mDERkMmOgTd6/675SJ48xEer25ydCU29+J1GBfq
ktkqOS/80GninOx8Yn8qhMJKLVH8BQplDb4XlbDkcCyD4k7m0n/q64vK3SYdqX3/WS6QYT/bFW+0
2e37ELnqU2uuA+v0m1e5yVruGePTfrndd71110YgC15HFnRfyZQcFpn2wAUm9rvAUG6VqipbY1PW
vUCKiJdcvd9I3rwR3B990zQTmQ14Y0K/e0lc/PQ+S7TUUFGX6295sV8DisZyCS1EpNgJmqWgTs90
Kwi36i4z26OxLwA2cD+vr6LAtkn5v9dQn0EPmAvO+WOyCnxprCWPjjsmhUtITXri4uVjrMkvQ5u+
zFJXaExqlrRYD2Wqyr9am6G6jGrKVz6Z7hPdUaD5icLCT7Uqly5nYqr3d3EH3lWHbYrnFQuGWbLi
pmSmAAZ0FYMJPjl/CCVwnYMG8q7en+kS9S/m9PaRJPRk7yXw9m2Y955gIaZDVG/S+PP2K6iuGndg
ljbm+c3BduB5shVZmKdbmHskKFsHZMUmW93idHrLdIY8zsjLj92rYgHJbMx5b8h04s8gCzsNruwR
sr6DS2GPqazYo/GJWNrM7Nh5ElQwSzXu/f4P/67o9FBJeOAq5N7mvqgyiF91y6F6c3rEQaqmQNlr
kV8nDMxqnBRx0yK5blbkJORG+p+I+N13kz/fQbhUPOvx2sPFRE55vhnYyiOFz5ymgEIANohaUvHJ
zK0VChtvDt42fy9nRL2zuRld3G2hhsEXqMN9fVB653fjwxUl1SC3b8sHfLKQf30Bdfb+xKPVuCWH
lyM5BmNtYH5DUalQnkkBoU/avfa65IoGUsRRotouptA7Ga7hqp+EsHvZGnZDC/qWKCzhxPKt3ISX
tgeguI2CjlDaIUteNvgsU+qgAa1/FIzxcUp9koIU+WI56WcY4Or3QByMk3nHxbHRFK5+n1/XFC8A
Pm83pC/WNQEtUAJrcLutJOZmDZ7fH7cqG+6ticWoTd/69Kvc2whBIMi1lL7J0pXuWwvWj3K3UdJ8
0si/vg6PKeOc/L8QYq5xmHnZLkpEXc805nSEM2UsHGd5KBnDjc8r5t+rG2udrCKDJNnQyM8AhJH4
y27VA8n+hBBjwcMVDMR4qGGDpwqcwHREDz/YGfk74CqxnYLkgFRxW3NMryYfNB+XREa3WxKRL7Rl
rnE91TUT0Bfbyz8/j7SOhM9C6f2zHw74KMB1Btu/VhSdvKMImfalSZUL9QclMQwFN3UejPAt8Pir
0CFHhLTcKhqCegOraFRceTqZ62zAaCNn3ZnpCqkapnIJVFzzviS0Xwo/7o1ZFeOt3g140uaeKRHm
LWyd4utWqG3xJ1S4hAtUntt7wDNmtcUG7mKf2T8xW3dZwA9P6BpJ+XVH0fvMuCXj7qr3Kkb9UCFW
HALBE5MAoEQH6gu8rrDihC7DyrLdZ6C7zG6FKK7a+3hstukBCB65uygtidytt5eiCA1hIW7FSfgJ
oD7qqOcFLKUl23ysmLt7enBzdI9mj5218J0wCWSuPEJ8TQpZ3GvfpEKpGHECO7aWM4YmFk4J6LUF
6cMsLSKuYARTU32eTALk5f0Znuc8txxGuqLpAzgoPnJviRTmpkOsoQr9sLL6gvdjMfExsJPvL57F
CPBno51hwIVNuipkCOO0s1LXqX6JFvTrYrrztNwgc+tLEbTvWZmhyCYfvLSiefLz7qAPigtSaraF
3eo+f/x0YZeoyx3kbQeTmAXJkyh8U73NMZx2vG9NeY2iakR5KgInB7Hk8T6dCdW/hcUICBY6hp8h
YEzS98WJewioU9/a6LuDo7QeCH6nFDNERee0d5f3wMxQM8n/4/f5hiForKEpJu4tBO7aqeGalPrM
0hR3E9K7U6BQHkgc4+CJD6Bic6QsfvKDa90lXClb/2UjmFepo4dOxOzgfA+0CSSu5mDV2gD4dvfB
LMRYcZGtuc3Gu3gJPV+Ncfu0ftxPg0281LradoCcRJGKz4ZkbOndWXy3HMJVQfSV1egIPo0y9B2N
xv/O76LNjb3kO+oJncsZpr8goMPZyaO7cqpbtZwQtrFpe87kvcc1a/+PsZqzJGWEUwGTRgwbVyh2
l9CfkAtDOMR3IledKKTj7VPF1zhMVI4G4N0AXhkvp48wnJwWqzCI5Y2DPuR8xPoJv1oZdMmM+9gP
kPzjEFVuuoBtNvys00Rd712V3iX9X+cXmiT+o9y3MSt9kaI2u9kIxH+75KMhdwIXLMXTSYXqZCd7
HvecLel1CYMG1oNfEUO5nCwP9XzXy1YUuzXVW38D/+Y35ZDXdhO1mspOny8xfZV5HQS9QIhVJerQ
fjh3SQfYpf9File9a5Cm7fRtces+X9lQKk9YH4GAS3yweQNJ4i6HUdB5N0REixSRt3DlUb2RQePY
kP3QaYsii0b2XZag+Fx1EkvzBMxxxuoSi7he44+47TfIzk4qdGTxxjUWM4HVOK520tKTtSNE7sUN
PcWlHGcQbbb8OzVW3IlUDcQxLUHWu2ymGOkqRyIWkGJtBzevdU4IY6cooXGYlu1epBjJOEfpBZyV
YJpLVfHHOuob25aFNMHrtNLAbNTvpAF6VVa13jEDO5rI70nXnwfYirfJ6Rtwh5HaJZXAtbZpue6I
kYkDqh9lQKI3omwqs7anA+KzxxqGO6C0y3G1xkffBhWK/Dyhd5Hpod/sSz/bxyhoAXJBeEIibz71
xNc2JC9HBjod8z2cfEdIAIfrb8tqL9my76bqJbUnCh3lXnQ6x9SsxOUhsVAmVMeX26I0vOIAr11n
/J6L7EhdGxZq17Pc2w5fxuDrd1K3loe8XH5wx4qRQhAYKs/AXmiyoVK12FlTjczZINAWefOEEXUc
mvyVOHKUi34qihdfISfhyz9P3hy6RmqSSV6SNtEeMXzXKDIDkjlUzVrcUunIWbjWblhYgfRWsW8u
IX//jt7vbefH7G/CYjvb9tYO+I+gHs+WD8c6EnK1WtqG1APYKG3O+ByyPRt8e0f/ZzlkNaXEoKw9
FN40ljQfPg9pl81XPbTxLo4sl/oySu07SZ7dQEtASfv8GQSq9lefNJnTacy5vVi56Ew+VlCn/tF2
fQzPNae4czx2TmK91BEuf/Wjd/c3nbptxyQUhfrbBmpeP2yCzABps5CydzXTm0KacYOYnDMwMeXR
cSI5xnxB+y0CorRPX+5B5BribQIcszo8sVpMf+v74e1Yg0VX/am1HoauIzDGDBWsmbi9Ir5E1dvW
kWLYMXARVopZeml0qrTCWdyGU3FzK0JQnsPVB1CAXlqh+8jT2TspQ3onzU5yaUm6/AdAXsxOpEKz
PqOT7d/FnMgfMhTaPPb+bf+V1QpOn9sePfWUNpT5InxX9nVucmQujbiy/fG6qlh4QkU2RUpMmCIP
ONHP2ccSXZoveYlZSb7CWcITYTbDZgovk2iKrMPLJsURm2wn1XXt/x+SM8th+2+lvFfyvNcfA4Nu
qbFtQyoCKuYYrwEgr8g0Vgmuc2gCuDpODChQL7JjLXUKbxdSzLPksX0EV8kHYlpTkwexw/6JRxyz
6UuuZceV7xKKgN8CGJFSCz98sZJpvOTqefU3FG5Ic6p83ZT6mDugUsUBUhrZrTcoS1NPWd7s8k1s
I9GjFTvt00iPzS+OZMVKJpWBhrAdSxNR53x2iW+vSyEjm4kigfdc47Z/zrJqYSot3Dd/GGOqkgtC
WDMK/HOXV8caQe+b515mb9cXE6Jk3Pt/TTj9d90fMmPeQq2VtS9p2QxZEwu5T+lO8QVyHqUA7Gk/
oDjjZuN8swtJJMEtUA/bvlxxHRHVPM7M2rPwDZl0Ql2QgnnEM9OTSztUvVPqnjkWeMbmCEbDbdS7
2zBT+aqlkvn93/qunpDob9gRijwsn7jMuIpsgCjQ1nRnhHK4HLA0puOwxoVZaVHqALneIOJCq9jN
GHelwt+2cWM60oMrPWRW9GO9Alk6SYNL050lfQ12ImcrXP7MkgKUQqEoqVFvt6i2lHg+Ud2ZlTSO
stQkvObg9hK6Gf2sIGHWGy2NH6OR+vqA97eXGtXYQ+WVH0lY6n5Da+ujsPptp5vBEYW/d5Y+KaOs
Bcn+1gppc0qiFtua1FA+tlGElYlXobOcbtCQHXIQwjjI8vo4f9rnFV2Ffy6Hs16gx48uZEyzRYH9
dHI2Mp4R1b5+aqdkPyE1pq0uFaZX+kucGnlfTr6Rn+PXibG9TWLIhVwzEpZvjcKO3sw1IgdiBH58
5Nr2CYtAJjxF3UAKxsVSOiUfn4nfgv1xvB7hcrBgwNJcYrx8RgzyiClZ/qDb5ca97XFIRR3aNUuJ
tknNrafsMM1DwU2SBrOVZE8W74gARuGu5Q7jsnUVTAgloYcTcjJAp9JfdWmG2K9tZtj4sWI94U5Q
l6gs/Ys0MdeNmSY8pBJgZ0F49p5vH+PCYHhrIa7PfvLzDmJXGsflbsJYcRLafjM99WPRuYV5EULT
nmohzLSyNWmRoSu2eiozMNiTngWCtNXv+9JdCuoVbJ0tj07JO06GPNO9WirHFq9g6YolerrsZg/I
kQI1aEnjVehNwHBZVmWk1NcW2/j6c0DLalP+z954tm8AcyQ6bhyFqPPp3sRGNANy32YDe1TwSdXk
pTYqVEq9h3dHk5a42BfDGqapT48HnSDCb8ly7Duhjgugje/Dwg4WRPwtcEnx19VNHExWA/VyaVQf
3XEky7JBD+b9dU2DwMACAWsr8Gi9XQTaruRruJ0BVZNmyJ1RmGa6LgCLg0juZxwrwYGgMKwa//z4
m5d4nbJi/6EK6XVSjhtzZjMLFZschq/N6isxDXDEcTyoOtQ4hrMkU5OK9osGXMd+jklKGKJv1xHw
KapvpGyRhp3PIuUZj3nndWP/btQmIK+PLSBsIHQ01X5LUJSd4NwsUDm+G2bVUHo/93NcYeNEjZLH
BW6I2pxWdHYB7zouttPa/ZIgHwFgNQLqRZ99fP0ZBGJ6x4wFgmgb3YNFBYPiab6wVkGyotcl/jXf
caPBKSPmy+VTQfjwiFSYxzqSbycvgi+1jrN4hjEvWc/n1dh3ph4W9FHlU4CFVD8rGSpFb+BHw2JN
xlKbdQIzXuPt6Mw21/4CYa41jbSezYCmfarYAXULDNevhxw6U3XZbIOsJX+2PJBknx3FlCJSqI4b
W8+cuLBnnoPM1DzcEo35kHH8wGDUJuw2daO+Wako0h4D4iWTdNd3tybarsbMI/X74fwcH2gm3bHM
MN87r0ybN64AF5OGgiinO6mfoMJBnljP+ovx0LwCAR6oVP2OmuI+n1+7kHwD+XvsoHzz8EAAZToL
M97UFywENe00O5QgZiNcaVi6N1yTpj2PXftgS96r9I7KWCfOOZvrIzuHG/v06Jx233N7fEMgMtoj
eywiMT6rzacS9v2MHua+5+XZVVk+3wpO8bi4pn2zP5nJn5ZBuYFMGI/kH+vVkAdptQPd2zh/mYh/
o3RJoiDTzXPz5tZFkZ0CD/03in638M4UYwz0cQbr1ICJs3E/Ab4vq5jzM7yCmZfc01tnusHbQ/nY
I51eKfALgbviTMrCU7AQdh7grhY8OOJqv0ZPBCn7W0sjXVloCkN8KyoicaXqOQzBrhikq4sz1xsF
bQLpCwkcGkh9vEKRanFmhB7GMBZlRB53ZFu9zB3RKrrebhYQwYgNULkukCatwan1bYQVjxrmoLDS
dGDhecb8UATprIjFnd4XOMSwISlcILKdF3jaCs+TiiU0fbWGCaNO9qAFqfuRv0+pCR1y5khBAzF5
X3SoP/QLOOVJudfyoVOXwm1j0Ol29VwxkdlFrbd5TV3nY6qycsp3DGO5FWcdEsw4jSXwE/jZ8OAH
fC1SXXZcA+umuHfWn8aUKMlhxoVm0/2XvbX6ZTIg4r6wtrk7AQkUUO2eU7dcAJSUAuTWWywd/ikh
KC9DP88cGT0lXsdtEBv+rWBZknKBt4TFhxiBYv5/7SwXS+m0PuQiUaHSXbHFb99sImzoz/gpfT0G
kJRhd4J8OAB+aVQ4dx0RGAeK/LuXM/2KJRuVXAZSRambpWVsTDk0rtPdSuMyyKaPX+ae7B7WyqeX
ArN8l5rL4FwIHrp9j7m7DvCkAygJigFmwO46QRSUMVbzw5nVRtyzp04myKH4tnx5upK7s6tOjDFK
1fK+c/Zw59mIsGnZ7UHT4AqL6XDpwD8igbVOKeYow5tE9bnlKGuwd6pEMHaFwfY2pYyle7tfWuw5
Yap56AwzcT3HMXmwRPPwUOqm8syZGwt6kcWoRGVg9JLFBADcPbyVf7KSvz3oYNVmgzNYpXBRSziU
hzv368isQ/DVpJ0hiRyU0/IOIrflZzbgZrWoMd2D6TLNeJpkc8XXpcZkFZccECSmnfi7HVOzDzI3
0nKqvThFy0BRvqNXBuKFsMW4/szbuRXfggf8CGWHTw52fj/61HepbZD4lMrdSbgX3jkRVCboI0Og
bohVWV/0CmFzX9j7QtInbGdeZYRv5KtSlEdKAT1gUlJ9TRnBgYD5OuVSc49ptJqkByq/UodQfkSK
OqHyPHTBvBdCSQpUbwlkbRY0X22CHCst9SZh+wFRzPBet0oeRPO6JdvW0uWneLORf0bTFZSqIScR
ujLxY1awui2uc0mLcOe2BwVbS3l+r6mUsHPgrL5AzGSU+1xuKm2i8gP1OhK4B1P42ZNwcHnmR2+h
LukqUwLwZ2/MiH7GKZXsfTZ/+13yV0zjMdnl2uk7eqg1KVBN3dqpkTggeoB2njW1m6PDv2ODIqCx
6Qn3LOCr7flDaVD57N+uurex7UDfW4QcctRv5A0afbVQGRrlJMxXFBQ63fSpBmQUyuDdSNidyYhk
oHgEeI/SK4HIKbkA1Kiz+NZKvsfjcAzRFiVPSFQsR7yzwAPKuRu9RHLHfQSHuA6pvRGaMD3N2fG+
X6XQQIu1A523zGRFbXIttvdxzNGTcEiA15/IIzfpJMLj3AHzztC+q7iJ4H+dSMVfrqufZA1s1ZCb
epFznwUBBX/aL4mtWZtDqnpxjuxRmNOumwwLehxpgOJ7wmk+nwNvSwbwOHD+q5qNzcZL3JQNpFKD
vIREL1AJdsBiKRXNj49fw/j/nSovD9dLxSMF3bQmscdiKJulQRe6aDETutIPmfpKCLSBAEUZjRzj
B/H2tnlq1lRtv/we3ZWWG1UBT8wrUKBqYnThq3gCMGP198MTEnbTwG6jNFzoyPRdx3yQYVU/fKiF
3eZrMSWlD5k6vqLyUs1Th3s4GCAAFFY6I1BMwIyB91p3E6UwX7hLWHe1b/zZQNOgBhPApHRuMCIV
U/iLytDaQPvOKqgoVNCiqSK/N2eMH739acUu1/RdxvNZILyE65Aqrc1H5wOdeOhYbfnm4jaGUY7r
jZ1nICKTmtSi5LT0Cg7iFLQj87zeBgokmdp5NJF/bR8K5KQALDkv5nv7i5iN1jNfulS5yDjO8A7/
huIAFOMl/tjVi+gckct9YvR8Qb3XRc2i0XBmsoc429ToQJZRQEyF5faeXVVHeWw0X3ctzpNdAZMf
0hmzw7ckqyBcNguW8KQA/8GsKZoi/o65nUxnJKc3Yr4q0z++PicZr860ZrS0La4HbfMC1LoOlcng
T2ZgcFugs2h2CMCBYXXrEb8bDxjEIZi0Ci9CWBb6V/TXUkg4SPUO90UWC3+Ktx+cqJDfITcQI3j3
wCFW0h+ymrdr/sCkf6idNU8w0+UQFbHZjBIRuQ73zXSQnhQmV4KhaF3V9TuAwSQQ+6kO8+8Gtuvh
DbMk4Q2agdfeLXK3fNgfO22G6ZKqEXigOWbKwuDG1M10fPBpyHXjRGnwD0IiGpLOUrr2RFQwjDU4
8xxhMiSn4zrhz6S9sNDvV+KHamdCEJs0XxqNzb61NkvJ2/Gv4pIsn/r4SlotLSfLW3SQZctGwg1A
T1d5vv5kaEs3wMGcA9XokJ4uEh3bXgRtn7WUuPZagbZBSq0zejI27lrHTgMM1NCL80kJTYrubZYY
ohNzTRSvFNX0Ud3kwkytK08qmLX8tebZmJfGX79r2YClCIvLSLxlFn7y0r+5F4a2oz9rdRRTExCU
ZuznSPchyNQu0J6LvpX+8lo6fMP1h4OquBTL2L+lnkfkYSTc/Uk8Gog8DOTmlXfBFxB0lf/fLOIZ
/Lqz051c+dah1b/w4OHs/QXbtMF0nCSNqLeSmQfkATwy4u6ehDKHugy5+/6KMkOUfRF8caOW/OBP
aCjHwOoPrT/s8m1mGKrpYGr4Y0WMvotZzDZw7a/NPtdiajagy3njGT8IJ7t34UGs0oW57+zYSRU1
4E5MSEqS9nLbywC/Ztwvtkf0+VG0j3MUn8wZDFUAbuWqGGlGF/TS0Pzgb042ZGM4OvxN2CVVt6SB
Q93I+tGN5VnBRhypQ1Sfjecc4EiIi4bJd5dYbOLW5E0W1qq0TRVfjSRip1+D0sVGFde0elLaiCgd
IcI7/nDDBDQlFux/+jSUaP9TFFS/R2z6ZsxT80QYcxtvvAN1YYCJFi9RT2P5FIZQVWZVAyOUK9Ed
pgYC7rDKWFemBuoAUVopO5h6fstZeUvecXH4xrnROXaWp5P8iRi2XQFo0KE5glK8Iy8gzvhvljki
aMARPo+nl0l7G17h1fqEJZJg60504hp24chjpip7Bu6FESSUnV/IiFNfLu3+0Pt1yH5R9uJ02cD/
9SOc487WVXAla8EVxuBOJC8m7ruMqAHDc4JlWkZMkRmCfjGX8aU0CeQKTi3NUorKc8Z9RfF0wOjL
xWc1+Z4Bw8AL3SIEB4N4QkHjN3Y6umdH/b4hFtrt/cA7NmuSzNrUTEL95BPDyS9dt29JorYNS4iE
Uz66HJhTmGW4b18m12EHiBLMEaoen+qAP3I5VKJOWeY3DvDtXm+yEExyeNRj45tB2yY2M6N1yg4u
X7m1N7ntapE/w+MpVDhtTVdT6gH9/MxGdxl2gHzymbKxa0/YjVbOIxJLOoXbes1jLDH5r5m7TPRF
ePiqPaDyd1AEr3k6VAAXlh+c+q9kolsosqZIZuvQW66LkpOIQ5Mp0BoA4OoBzuozYBvyWWiQbSin
Oqneqrv89ZsKnVbjbH3Q/dxe6TAD6HxIQvfJ6uS6PGPCwgWKzxqVE7RLJtp7fWqizcXDcOqZyr9B
PbWAM3aFor8sNb2LhTPr3tapTDTz73l1kfmWZIwKWG/ovuYl4IuSURt5Y7IVL0lOwgLiZehbn53d
zROYZKSfbnKQkzjDmTOeYtbbbmoF3iqIEjY0ZLXlFZCpa4/HvMqlo2okUd5o7P0FTFQPWURTg9GE
Ce+mfOVNOrM3eiimrMQtl3XrAqL2RSnz0AhA0sotedG2WntFTNUx6J7KLcZFVkGgc5lZ/F1tl159
6vSStSD3RR+axscOKuqT0Onty9wVfvEwFyjFvCB616CohpaxdF9FMbWW0BmrmV56iLXMxp5ORzEJ
9YrttgRl03Z04YnAjGNfulA8pDHOu6g6oodDbLrxibtr7LiAS/xn8OfE6F0Ye/ydMzVYbCdsR7tp
nqNm1IqDGuq0iD1MlDbc4iEtrs7E3Z7k58PRyjgNXlyTTh5YOlXQCEqEBabTn1HVkKis44C3lY/E
LzO7Ci4Ququt+i/cogBvByJutNd+X+3EFvcxOG7motpFYZn2VWA0chvT9Litak8AFAnSISrbrDOq
l0yN8p66WKlLBQlBz9IqNCF85HsmxTC+AWpD5F/ub3eEKfTvKPMmG8R14BiOlqjulgUFSMjIMDjC
VesrLs0yDuTRC6bgN+0hY1LIK29y3nzu/1R4QJAZpqZnsFVKPh4aTdf+TzqmudmyNJrEjQXHyoJM
rHcWI/dxvls0cTgs3ng1CbVk07ay1sSSbpV1TgyJzaovO06NgTmct1QmGlpj5j85foTsMkIQtvjL
Mzw1gH+u153HHw1oK4u2+dQ3/AEFT+kP8iXQLu1/Me8IHcuCYZMIH06lC4xoVPkCTi5Z531+GeuM
TL2zGc0Aa7PGmdq6tPSWFZrlYQuerV00zJAQAXUqbQXCS+pzXRKacwy29in7wSrUl7a+QGPU8cE5
hEIYQ9k15iL/Dd88bbG9OmK6aamTwzT5BVHS/6Kty+uyF19KbTmZJM0sHUd7qWNCOhn7VCOLLNDQ
+dMEwePVxvK4oUqTG1toGJ7TlM52/xrdqNXet7YZSgA7iG8+mwPbO43q+rzjgkSGcPPxg/gz5h56
jFSad+rF3bwPLjmy0+pKlDaxVAqVt9QuFiNxNdhDyy38PjqSRxeLVFBZjfUnnzZsGzTDlXfac9iG
wb/1wDFGJUVm/cv+pkEDRKluYyBpiMd7FTWaamUPxt7vxMpvYtPQ7AgWaVv+7hZ9hCCQColZraq1
R0wFIE6bntIhuL2BamynS4fvGJHjlZfFg9R6n878zDEzw3Otr1OEsW6e9sh78PKsnedQ780BFp63
Ne8zhRbOMccT/dDOewhMteagX1wim6U5fNzrl0+2sUltvQtpgXiHh0XSV2a56G39E9qeGXZDVAW9
9HwC9W4Zw1hEsUX7eBRUgugaFpPQCA/MxZ883cIYgJGz0BzvuJGFrCJcyNXe82I3Rm58ho0+tb+4
J58MVkuEOnGrxPOlnVamFR2uT8fA3hkvou8RJJ+YxdKatxo4sHzxDkx/v0bufWLH5jjjyoCc/2dH
TpgP3VoCawqY+F7aFwxebugbKjpXEI2+VZdG7/HMSCVJ+NKWH4a0Ixk/rK0xaklIYo5mIHBGSc4U
zdRBAImlfbWj5/Z8phImTr826kjMaAh4ivo0WmpJKXF2mtVikN0xfOVj/1QSJ8AQOF1oVg/N4cs0
QV+CaVpJBjgLH+BXIqLZXgm8XRWeivM5fxBauYos+/4CWMih1aNn49FmXtjxBejs798KwtngJMei
9Pa7aopLmDQTNFKxc4RA9BJnyzAnM8DNopgIxFuKBWRLrliEFYs+xXPAjPHYL6xKZetgHtr0nGXt
LXMyg3sLOQQWxmbyI09IGDb/huNFw3J69LMC3ghR5CTyBAVXTu8RXzTlHb4lu+Ye4rEKCDrqetGr
fd0Nvye6uagwfkKcWWNpm5Jon+PHVRt1JuDlZqsYaQcwm4AkcEgf2gO8Xcqnt+f1j2V1rcMvBO8C
Fo+huEwtPVp+47CVbPcxufEcEfQj3WBTIsh8bpCMtVjuTHmBN5whc+B7L7dAp0rJwQ2hZ1+CFkzb
NFcxMl/7Hsz3j41vaHFxifkfQZIl6DelNopwiTMvzbMxSAwrymovjDWLQv6aZ3CPcjUj/txjkYVN
2cGMHj4WjgCdvuGw8MbjYTPIX1fnOuhBXTehHsIQFqpABRcSanr7EDSAs83ITx/XProg6OHg6CTl
IqB758m+vj/PDhH2YxEjJXc4uQo4sh69BrCMQLNiFIuco9Z44l/W6c2S5ak4oyN1zqADsn06WmZq
tpes9yBFVSkuaYuz/cbTO89Uw0EXtc83KPmU9Xzoa8meAOm4LRDt4/2L4YqUqE2xbtD9yj9G8WR3
vrFjnMmAQ722EwByfMRpx/DRLvM2DxbYGoihM8OioI5mhElMMVcjyVgGQFrIQRvBV2SNNHY9vvBc
f8qYeJmhIDNBUKIGUdCR4uutWiC3SwqMojH1JGSgNtX2aCjDBHbkSkKgUKmmJBK36mXgtj9RI4S4
kex9RVODAhggZAHS9g4QGD2tjWSUr/NhU5Hdsr4Q2Nn9gSd9DqQzB+X8GfP4vzJnofshZR+qzda3
T1K2GAhmoGwuqvLJS1PRI32eovmIji9R0KjzmqYN9bN8XjXmLzPgsOGTh7ZG6SgEo/2VB526eaI+
NU9hdjoCv3aqPgn9/9lqy7uwJM/9Prze8dATbwxzEbCt15e8VVmNG8HZnGAYZ3lTY5k1Lsx2wlJ3
DXyPkIyQvuDwL2u0V4sohC/DCj8oZoSKTXOt31S/2jckchu8fn4gyuNLWQYQqJyeViLbEwjE4dqE
g4TBxeQII7BUnIykhLtTslYdnZzq3hlSydOTohI9vwR/R8kGzggVy8enyq//++FA44n87kP0tzFb
f5FrsqXloeaqFhqbZWB7Go1yPJmDpcekvd4dNZ4JVsLn4p2a2UkdVbFYFI1ZJSE6mhXAJNPYzDbn
1a1Jc1x8OOo638yIInzs7LDCcnpwO3QVTsB0ZWWmKn8HgejYlThVbpAbrHWZr8aQLnUda/kCdeml
EskiawhKLNyJF+XYLw0hjSMzoq5Ig7RjWyez143elxtoZkvm2vgHImiDs6+vB03/7MXYNkEZwmQ0
07faq6dYcX7Bio7MzlQsEMIUJ9hKmCnkheZvCtvM1twHrDGzlP6MvV4b3sdBxUwAkGOksbZQNHBR
FUMG+4DH1ZiOLGuJGAOrY3P1e1VQaz7io/L3ZjxF26K1oWuST8vDbcuNfzz0Vqc3mCM+1vzXOCl7
6iGD/NVKjMhReQ3EnicGegMC8YcUYsXs0trKWBJslfJt2ibK94S835LwJZs6sYvrGsZ7P5WBvz/T
1K6jLmJpVnBLeQRAnsNkfNFqG/pFiNIEraWgkfnQL3csZ/5lhck4CtD+QYeFjNAfBeLdA3faUeWL
1LY54VtlUHv46HBjn3MgFrEfSgTBEArM3kdJj7J40PvWTAuLkHGapvL8SoE9P86cRES7cN2n0GLw
8vTng5miv/8M2p6IS9v9ULTC2BKUoNhZErgtyqqHUiKs2XVL2uDvqUXOBBnUFMayn3odq0993u00
L/U1LyT449k5Kj3PT88lYoQFoNMm0lYP7l9EPtajyA6Cu7J6JYMASJIxVV8UN8PTRWnLgPrccuHv
OWNyIQcyP+Mb/e/ZactwAhBeWMkG0s78ebIurMxGKrYOYG4zuMfrY5LoTil6W+y+JCuRLx7yYZ+Z
w9s3zMPDLywtiChlveGtWrXby+wRpx/Be7w5Tb9ObWVN+KBiJG/52ysymYZjsfBSSCU3rdj5ROi4
A3+Gws8boQ5TX41fZ1+GtVJl9Da7e9YoUBJoSrk7s9RTzf2PscIsLUa8Vu4mFo0Vxvuh3wqHsM4p
9J1NTGM6Mzr/davVzA3VXSuBIz8NkUQ10tnhgOo+wgXEVqXyx/jILC5sIWdn7ZcUEGpSZQcL+Pgt
ny9A+bKlyII57qVgLqd0MylwAgo0vrq9pEXpkP2AtuATA/K4bEkO0SNQqKAThftdn8kIyWRD/rsk
14UP0AlDb1pCOvJLLV+8C3uSVJhoWksvKWc+SEh0fsA+EdwWeWcWDXavv9eIcQJTjSDQWr1J9V0i
avKBdgagp0hlG85gqFHdqP4ceftNAOiLZ55gktAZeIyyttu2fXNNtIrM8J9f0QDKrEtr6e65DfVG
LIbR1Vi/Oz7y82zGFR8V3qRc7+r1FH2i/pqOBrSbP5aG3xDCF0/s+7YiZVH37Mh65VF7XwY7c5rC
uvNq1EN5EIxRGKz/gY6PMtXCA6i4eMhTWetzIMRyj9AB7WkSjbxblWzDrBdgz/117/k17E3DXWta
zNcyHtvx6vMQ3AQ7icGymeAT/pBjAnwVATD+WfPbaulLZk6x87BfkMDi1Tp7qBUUOw1NWPFfeCz+
WPIjUEQUed4F1aR2K4vrPFj5EJ9qA5YsxlLA7Ew8bZjAnQTbk2tc6fRQZgfUW6V6nb38pF/eC/oU
V2+l5YkLgkwfI5dCPGSuTl/IuJWnBamq3uP3Zvi8GRYh62UXg4c61kPHmvfwFVNgCGISeL6RnOpE
ohCXyJGFTm142K9OGx0/l8Nkei4RK+tuDqMHLoReSqKNdA2E/+oKfna+9gw6ET+wzPjtCp/qjpNx
owFjI4ZwQhojaq9Idvvq2WDTc158xo5f6IlNuFrOiIn1MbBzAB+gulAFZXRDQtbGNUL8SINXN394
F0Pxg7iKCCStm0gpmjs5vd89FcT3kwjZ+hFwHKvmBw+V4T36Q5MVt4QuRKz7VGR0M86tq/x0EPVk
x0bNTb5p7jxvBsh2LMu7aO03FYSzINvu3ff9jJ44fszsrTDEA6LD8AExXcLqL8miLQKE6KJWYdvh
mueE54wtQL9ui0N4ngDq1RlXyywTL2Ix0fEnANCdJJdW8ImT0YIq0dLGSAWa3sa79x3E85+St5A5
YqKaXhVuqLH23dFoFp32wrQAm/jBqj3tbAJh0bLM0wDsOXOsZ8zyN2wrLx9HwLXRsylvZdLKXomv
QIVw1IAGmKnFCTtYn7UhYe0aBZi9rVNW+ojevSfpPIVS61Gs2vPsVdJIh6HvNdr/b1WYimQj353D
D6iBkHweRNwWGmjC8c2SZpRib8/zVmyMiTalxwSmed6QbN8zGYT54GJu811hnwunaaG6RXApGTfS
GcKf5uhVM7qahaMb5S87dkUKf8kX8rKjZ9CWqjkliq1m5LXjj5hbySRv3aJpoz4k9DkTTQkCLNYt
U5rWOSUnhiUMl44sZyNXCx2gKAD+IpWn9AW0Lwo6ItBJK9vTF118puSM3y0OfWcfDf6MwgjDe4U+
UW7mmRPMykkZD0CzltRy1hRyRuvhKFb2Wbqv0lBOkFgY3hqG8x2UMhBwa50iZppTpweZy7s4m9/5
QCPtlseU7h8aQkhzRo7j34TGljeI1KUKeJV6tYiFO9eCUTui+JLSMoGb3pZjZ9Q/1+f+vOgKTcrk
QyWXSGAwdsACgv+/SIcmqOAEvcMFFISCO1GqcLP31FzDhlaM2azskJg1AP8LiPCN1XMWctxT9URj
Jct0rsZ3w9xQr75aNZAicmHtaawsaBVLTaQXsG7yPJH9X0RBSzkMSv98zydri2nZeMS68PHUHkUM
Kvpv4SwramtbBcXqW3AtJHZ7LPHCd278ONwV2hylMWc5VuGo9X454AvgHIB7pL0TY8+cuQcute4b
JOQe/zxiQNdw4+8EyoJ3hh+BQWfnvdvEvkdxCFRBayx6e9tfuBq2ZUeLc4mm3cL0Fc02OSqJEGGk
Y2mLGKfpfn0Bkk0qTpwIoz7KfEAaW+NPFqj3NAiqui27CYEiZI/ylUNaATdjJScxoHvMgpf6bu5c
M5SU/K5sIRcvKJV1e9ABQ59mLY6nciHmCLf1qJonbTVN4migHKqPYpJvPywS1VuT103n/TOSFpO2
+xnZ2JtgYpLTSSzrggZx6xi+ySP9KTX+wnHk+LGt9QWB9KdaBqhtVle4IdYXYO7vhIiNUnz/hBny
yl//k6rQuQnmmKsyxoYD+PLOBHPad9iIZkzClAgSyIA/GM5kcd8KU7jH3pIyoZGHyxGH5olbM4EB
NqgpldpJrOCFe8ORkmUCymDuk1+RSAXin92aw3rSVLkG4vkjdE1cdtl+SZIIUbSI38ZOTEvl/qAb
JODu3pOL9tLImA3QsthgwiPhlxVEYmnDP8KLom5NPJFHUlm64OR65gtb0AxsYw1BuOduQacUfNrf
BZ/8nqKqPkdZmx22Ft2019j/HWukbGYjZc8nBr7Ef3/uFbXm9D/pbZIdcIZdzEjYpNDy7KgTzLPp
bqWdFHHg9c7ds2nnWH5RwyG4+dbelfZ+UYhM+d7Zv4K3zRP+cU28CkRZpKlNrkGlG3ikGaveDMdx
BmlZc/X9/Vy68xEo2xmMuOj/2dS0RcO8QKbDExbAaBJHik7joqygphllN1ZFEL9CexhcxAIIgrWM
7ZR8NBVRB76p6KabjVNOvN7cU5JMBsvmoW3PCXFztPgvi2FOgfzk2rpKU72jnugVzAVnWr5c5pL7
a1y5KPI82Ho15eMvRtgqpb6c+GoCEQD/DWIUKNmFXsnmMa9L84xfRsJ9rUXXsrwapEnvlcxT27BI
HlClr1mRU29mtm0pJTyFm8gRGXWLKhJvCfB22/ahjMIXe1qWjPW0RDbaN5KcKKf3Eso8wmjIxthB
2Wtv41SMjOsfFDpoCY2knL10Oyp0U1PrhVVF3ByvG9y0oMQgORt+uI6OmmJCn17VZgEjMP4/0S0x
cRIcuroKThePG+rw6a2D1o+TqxiaSu3Ju8rKJ4GVqfKEeeE+9Q3VZKkRbjl+HH2PlhpkIkfTBj1c
8mDj5lig1ZW3QldfOLaPtANTRCuz//ThUsU5THueb4L2uAykiuAkZdTEUKmc/AgPkbtz53//Nei+
wcP2a3D/lvTCh22tXJRcbX4i1ExSfkCxRELGdFSVc0LKRJF61rLEanjBHEzxipgeCmU6uczfH2Wp
VILOR2ZUgwHJVdH44v5TxZEf5T6X0CvNk+siaVstLhk+HkRKrEWOh98jsvGmpAgazbDF63tAd5yn
24y9JPf1hgB4ig0xJSNKxO1lbsHlhl/F+bOtXGyH3Ye592xL08WMQksXRHgZkVlHl5mY0/+4KqNt
USYmYrQ/xRGLXeTD5MP6MXN82YDueyQV0nIXH29kFq77YLe1rvXaX1Phmuulk2SGynsKHV7yTPUZ
AOZyOCnkyAonLalY5bjfP8lB+gQUEN5Jb5sY0juL/PRKsGvfHx7qSnY7a+eB4pBd8Y2KJfUFmlYA
qBlBFU21FATEt3jR/8HrrmvH1mdGdgxpw/fBpLX2b9HaiGc3lda0fJe0BUTqrFwD60p++GPIS3oG
9s+plRZcLYIZXFCPP4Xjt+2wSSdqVca9WmraAXE/nK+XpcT23bD6h9abyr0MWSXmaXJR7pkzti/n
51ikPwpAh4bRmCWuQPzTO+aRZzEPkJ5MHPQdNdf12dJlwwfjaky/ApuJVJX/mq3hJp7zl5glVyeX
EFngPXI+QRbC3GTISxL1/LtvIluBKe7iBJ/KyPUEgXt3RUhrJAprup3KDgQ7qEbbcgYHcEccD5Gb
YP2CCW/xD/0WH9b43nGgggFGsnO/iOynZWNBGU376lpfG6NIinEGHS7oFgxDhBD12tivf7WuNcyd
XC0IgFy+qrate/G7GRta7m/qp2/FIiFNndfxrNoVmJtOIos8t5FTI8BL6Di4wvwSm4mpIg7ICQ2x
NUjdsZS6tp2a82SXrseaFni4ruFvcTEB3Px7RI+bXXP8ayN95AN+2PRdP/2MxLToXsjlJV+ZBCr4
wplE7h4yzx3INr4rATZVVZyDiYX6afB5UfsRYQlt4AEx07XnorFHa4LD+vWHLOrlMKAgOUzpvoz4
PZJqhO+oiahNMTaEY7RJeDGjlzdi0Y3on5N7oH3n9Mgf8Rx+7y5abx0SDEh9AAO8iZfmYhpUUiYf
Mo9zmsRozex0dbbQyJu5b6mfiZqlaUfopYAVVw1xDiNG7tvC+UK2uh5wpgepL/sWNq78I1r+cIsC
BAk/KRZdpilSn+0f3sbHy880XUizPcUY01K9frnBiLgnIeDOgiI1lnYqIPG95TKBDyzZw17fXfQo
b7jysLcDA4eXjyyoXql45IrWahqX02ydnJu6YcnPBOXPQG5Rkn7cGWdfsJY+ETCpnD3PZTl7QtLZ
Pz9+kX7IsdimyUw3Kp7uiarYiYhZzfXv4b2N/0AbTx0Msl1x2mYdi1DgjGA0Z8dSZbM64ECVXEkE
I4QRkN4gLt1LtNHKV+1iIiYY66Jz629BKFGuA4YCmiH1LSIRXWMpgUjCTtGbwDAm9+qygmK7oefs
CiRIBtvJMM7YZTNpFk6Q9zWJiheZyG/FfMr9oNzx3Kw/QPCCUlP1nowC9ocvHLuSZFPvsGW7iis7
fofIWiKb6SGxOcN2mOP3QMtrXJg918g48rsu+uPjY7niI8x3yA70QW0o3PvZvlr2TOmAtWDjaRWZ
+Y/0/dMpvnhBO2EghCAsS6hb9nB9rr18yyz42pt8ggUYKPJVW/G2NOxGq0h6aHg4oikPWoJOBK0n
8jCHwkUrtd/SY3Z7Ubb6P1Kn3/wk6Buj35MwzRaPBM24q+fw4Kc6HifH/cpB/MYS7Zr0Jc17M9Ym
o0mS2tVRD6ryK+hf7KpEP7FX4XF2Yu3H9ZeD09acJ/zBzcaXnM3Uu19wNgDHbSEyxA1IgDgWTMZ5
7gVuOH0dTemdho92rf6am805KisQyxZjqjzryQ7303wv+YPtbjFFpNc4DQ0uBmJKVUB9Q2Z0YIDG
SC18uuOq8xef8IqOoCtt83GJAZWnZlnIdSsGEqTafgl/4UVLIDNiGp8NJYARrN+bls6o+0YoD/el
eJUIPJHWUGkQIuJK9W27MT+DU18m84jpxdMObFnwsLYgGArQMkOqpOWqZzINOwRnZGbOckoLjLPE
qOwhbI7Tz7D6dqLr2eKTvRH9TnliMtBn1y+EOEmdXtbI3LtB5dPmKYEU6Cu0mXRYr7h9hIYlyjGV
4mo+i/63snhobNj+ESXwpZ0ghlYmANKi8SlVGuRmVxmqUM64KbQyz/Y1gtIHvFAwBRPb4ElefQ3c
AlnlTmu50vvDyfs923O8Ti+FuHCNpSFIqLrBx1ZAtcen2HQ5Pa2FaENR8LaHOk6LEzcJwnpX+vz+
FySj1xJ4TKwFTPVpdRwa0lz3uoaV/EMwPviNsAA+8klbeh5y7bpyuXBgDiwFfrYMQV1Fb/FRrkmf
gNdLusB75p6G2YNynVJlzeElBHW90FBk3cZjfrWYaKV81tuPME6HUuvuuky1al/mQscld2lTeq+O
nngknfOh8HeNDL3KLySpsnAAYTSVIB7gmdr80NGJTjsH+HBT7pw+o+/gtHSHvm4Hr63PWoB5aplr
l9Ei+tRZl7ehDig4WW2GPlAyzWwHB6tbkUXIn3TR+kM3GZRwTG1mP98mnDX5t9xXKBfWu0XQvHmA
Ic1CtTxy1T9eCfNa051YCU78/Nxsti1xvWHAMrdPXfS4celq7DdpOXdvJlA9DyR8B3fS1ZhZHKqP
YMFu/Fy9WfSbSwJxIdIGvMcTM8fohJTzxdTxBulvF5Q375ZuQA9xb6R/BmKkQtSoQ/1vz79NG6MT
MTKZEy9Q+YSEHUWGu3SawUlH82FgoQsOABSd0iyGkL0n0Pu24mGg4ynLnPd79g6AdSswLmXdIxvy
1EmcVQ2665VgQkAHKrkIisloF3qlM53KN1cCZ00kKPbSB+Q6igwArQVE4C9kkmEAmfnX8UxT9xlK
cC55kuilR5KNQGMUObCLzR6el6eAHCRuQJP6TwQeSU5InI8aPy0HjXvs00iI6Ucz1djKMMdBsqQP
iSevoP0xd25XvstjB1hc4/kxN2rMo8x67wwTGDMuhRKLHK7hf1G6CbXPfuAa4OrhBmKId8sIOPbU
slsMNryjg1WTuz24FQYBsov8b9KWG3q6li4w0Dq74x9grFJ/y4SFGoN3PwzzVSyZo432NqZasuZW
ziKAyWVHS3Y9xO56VFsvu3pMvsIMdtx7fgtxkdKpK6t5weHKIYM73qKUzA++eTOiQIyqnBITSi+F
B8K+ts1fyizha4n/eO1Xk08JVdn+XpDO+S5hKEF1Hz3bn5vO4XUu2DPN7bDD99NX8h4aiTq2oO4q
xYX4SmgXsBikGfi3leVt9cQCJC9hL63oYJLsTE+OCdDZcv6wGsoiQRIeQkBMv+tQdzBmFI5kWtz7
ZPMxplTz+13GrcoWj5Y+FlKBCSHLP9mYpYwZUh37vK5vnjGMzFXcZAflVSGD2Erts3j/NNec/1ud
F4g9J5+KCmBZp4+BVOB1LpznO+THs/5jeP9MdDT3HkZdGk+FSv5uk7SpjslBz1d+qMOXTpzstjf2
ZAVVjWD4/QZuUgQkzagXeb9P6J4Jdd5ZICqKW1WUtu/1fEIIRmHH9CE24T1YskmpOqzQaEB0zwMS
l5kZUwP3uRwtVmYsOd+9ghVitg3HQ7L3Xr+rb06fjTePrAP9QcSCiQIBpLuFiW/hppgiwjfj2RWd
UuTLs7/UP7MXctaYjQR0Ivfo+ZsFY/y1Iblxk8vTi0kwMksZ6HX9W5ZOpzhxRRwfneiG8nNuRJnf
GwEvU3CE1BPUR1X1tIaudJACQ7PufzsDI5PtcxO6Baa4TTEIuscrCiojTbdhLFnFoRIiA8HM7tct
bW4kY9lGMWjWRR2ImcfEcHyjqZrNecsPaqlQWygJXc5I7UlCbCoO7nMc+iQIuuq0HL6YYqxkn+XC
+qQecc3po3rFqdscCfgHYpAW58+OlDHBMr/A0U2NukiOgeRtd8MJeLApmDRRk3kKNAuQcAlXld9A
24GjHcFVE/TnpIwPLDJ3tfnwwH+mtoz0lx+icBxYl3CKAKBvvxO6brtPA8UzeXYO/bLmDQj/we6e
rKzY6vvfqDNvrGfvOAkoklvtVfzKxP9ZHd1A9yUTrog3pvL6GxJ87Z9/TFiu2QUCpNsJ5gqe/s3c
hBjPFy3wy1hzGd40mM1u19wupzc0AP7aqmmfdB9cABEijRC1pX2Z6P3aALURsZsYvUxlzCaDptOp
1DfTqJuv3meSCndgZfd65RvADNrGuog39x/JjKbzNyOfbw3qK1GB0M539l8WJBR3cQeqU9xviC1f
AD8eq8oV5wvQgVcd0UnjstBI14YchIxgSO+elgc8NGU2CwzdeuL/jOeqgrNW/ZNGnMzWF+12lZ25
ATTQBjxsokxR7CUf3NaFLvBZCxu3WeWH4JB6tsa3Df0TQ43+qMaxw0UbGKV2ss+nEZkRyqMO00Li
bBRODl6OUUYlT8ZymNTxdmTnBCKEoD98YE26+ymIdPuiHjP4yq/AidKazuSW+/7/MD5BYug9Zh+b
WPOydbQ4EbUACFShadXUELFLt3c+b19mrkzIgi/Ku7Eu3oxOJ/hHI1/+xxm54eGR3PHTsOtPawhb
IsTaL4j3SJwYfewofyxBoBQ9P5CnHqLv/W8bEwjsVg3j3GM71kO68W0472eSsJH8WZCQUckyZ8sO
RvhqRmOEYgbLlBPpujy8FMQduDuBSpk8YV0llPDdL9kSJS73LYvXRtb8jIa8MFhZL3HHn1x0hYRo
LK1EGc9JTNsx5ackCn1ssIycEq51h9BvD+S7h69HJNYSnWTcZP9mBe//u8DEH1mtok0FkBM/UdHG
HMeV8KSpy5mV4e/dKbWXP2l16eQ8+8tF2w5kJv0ojNQjSmvFqZ1z1HEXEQTbY/FDLHzHP3xO7tc3
VE3uHYc7Nnx1NTV3DBppMCluIfcPRFaRhMg09QiCY2xh/DvCBtCsauJIp+PJbLDKm+JuqNrX4LvJ
IqzlRSIcufLwSsInA/NEf9nW/zR5CHn/3INrjpmzaxuv9uxldwzkhaF04VZpams4ncosLJp+EkVv
GEaERXn3BghW7yVscG7FBu2QdNFtJVczTruJbX3NzLXLovKlzOjA5pXjHoq5NJDpGr1Sie2JMyOj
7K3GwGO0eXUo+PwcXWEwn5xAB6MAQKiygPspi8out57krhiIf27b+CHffPh8vBMRClkUcCmlqoo3
DFg3kx51tTrZJ5clU4INEw6NvYUeXU/bsxb5nYRZ2coSSLPVQUEpWuTER4Cgjd997x3P8d3HGzFV
1HzARLjiqimu/AO30w0IenPSfoFispPWNVJtVvb0GbYMJyCtHq95///6NdE3bF+juaHLKOxk0uUj
GhLZwgOQtEHnPPIcd9Hn/nAA525TO5JiMfmv3Aqmm30Kzzws7OBuMVLx5sjTLo+B48Aar1wpOgsq
Rn8VNuXSjoIrIVSEpK4yTjm149vak0e+VYqrVJqAwHl6JTvRmJIEstsCpxnZNOWIY1VYdvjsRRVJ
w2llWyJiuX42+xZsneyXreBkv3OFwKqh7LtDPzdyZGE08Fvovf4qjWBmwjxwaQBUJZDG6dCOe4iR
SA3zwC/D886Zah5I7L5uSTv6hHNeNHaMePCu5IVg2NzadazLxs9Y5ILzSerJCFfdoatN1KpIq+uU
N8CQAOptZpnvSkDqCaZstyoBgGvd3KN5CabD+m9FpGRgaQqoAJ8Y7tEzw+tgdCbPwm/MHnkjvyg0
LnmXNhre0GGb89maW26+PaNz/AbCfNMyB98cDqB1IGg4+KtV7k/0W8apRAXZZi39JmppBvFwusWM
9CUdLQ76+frS8v8n5s3bT86BxepV9XhO2oAyzYkuf5ghq4yXnMDDh+5H5FfAh/WLqRysqA55VF4R
mAZI1nbL8H+e4w89DMuSGgnARQYHdLITLfwUqdHvD54UwBKtuLSkusMOlD+kiK0FRwX9z25CovoX
dvoocQrdq9lQniTDXW+THWu2OVf3JoRSELB8CwQqSFX8pq3Bche4KeqH6M6INVlzxCaiI5NxkIdA
TuDCrsSba5tA4ckeowsP5XQlyRrnW7XBxPRHHc/mk4zCiWxUPEKkhtOTCsSuyVx/3Tr0nPyNTYZ9
/7s2n1rJwqlnikp2BJec3NyWCW8X1TMS1wFt7yE5IQtAkRSa5me1V7IceUdXJxc0tXvVw8CnHj5+
yBFmOqQlhtHM9ldEr7Gl2mC2j9G9QlM4nnt/QQHAyDee1EyZZUV8ldR7+j0m0xSzFMIFV1qU282o
jzeYXw8wl2L0H53XYj0gjr+oSEOZ7a8S5FkoH+pdYR7XCg7SAc21Ffd7RpkpxbJHZUOGqUbZpRFP
75c4kz7hP7O5uMGUJLpVkMxzbMDkudtBbhUIpkF4PwX1m+4fAmtxCGffKXqgcrD9n+uCsFnyYo/p
f0EqCVUbFP1UDt/Y4YtgKQSw41CTZtBS1mG5RPiPVI7zp3osgR4gOPtgal3LDsm+ypnOJoXJ6bgI
cHLUFVqM5geS11FdoUqBpmtzU/Ynpl4YfVMTeofwh3w1VXXAk1ZSAeP1fav2BsnWbVFS2b9RvTOK
MxikUKDDsQXf+ldZAmgG47AJH97DQOtj2L+IukHPjg5FXgX5yRMq745mwLMjS8IBZrHfWBQEl6CQ
SlISpeGXVSUXi1QYg77xpk4mFMzCCZBKSzIj+2znKII+Mb5yraOu9C5M1chUwhD1WVV9Lm/V1KZM
F1B2NWQXlYCZo4Y3bR6jAVtImE7wxPPTpkt5Z9ZUwQsPloZVX0uEBb2i2YlfMQObMhj4wKE4G5/G
9nsKrCkdJycBqmzVWvwIw6HDUJ7qNiJi7Sgbn02XVu11mxO+WQ14dqKURMjPptx2aLbTQEpTEFzl
4m57i7BkAdF48rh22RMMyJ0d+B0DauvYGtR4OjhvFed7tKZw5gxOYDrYuDf7d4z4hFFwserSaX/A
23BMwtfSCoQG3VdOJynyLAL9/Pisf4oBYKIwLvClTb6Axo6Vrz0THem/Qr5xet1MBw1fP1aiZp6J
MKC2CdybM7m7pZD2dfqJVOvp3ClK/lixhvDaYdQNvxFgIPcpXL9ND4yHnwvhO829HFcC5LB6msGN
iaX+lbBQht9PezSK/wTtUps4gveiTtPo6ep03ZKU9XzCbI9VHfa1581uzPQ7GHIPtT4NnYTbnIlo
aDmKl27vHRBOJoz0LBuw/GDrQL0PQNl4ZLtTQ92GExu6djhvONufub/V8SKVsdbkoAh6d0bom5q4
EFmDckpvE//hx9St+f4+Ckq3GWIRCSiQQJOM/BNou7dUWST+VjxrOClnn4wvk+POerxCSlmynlKO
g1Px19ElEPmvDyIfw6uNZesaX/RQ/IUgak5JOEzMtCIDKzJyCPEMwDSQup0eaH0ZZ2w7A/8gusTi
GkMus/tUEQjHYINiNUz82Kd3eGeu47GlA0zKWRBY5XqWAIuqnLE0TuKRbu+2l3JjImivjkAjrUnf
yEVtDziGnsObX0Xn654Zug0+ohZ05AG6YgbjDugj0SxXW3GalfLNoOHlYA8DOeLkjM1eKMmaWmpt
2Y8hBeh5+cbgqPuLYlumpdlPzbf2Va9dee12pkdQDHDNfOlqG4qUMS+kew9WNxvXZ09yZaCSdZNE
0eeYgkm4Wm1xQ7AKSUTtyw20K6kaaz8yJactYMGj80K+uahB0iC/Sx6M0fsO9fuzj1Bwpg1GFM31
DYwY+frt3rmbOLjmNND4z8eGRwQW7KecWNu83w7LzfrEuCTCTPwL+vvAS/S/xZll1ojC2RY3pcOm
YLPxNbNcgRrgde0s0UBDYEOe2M5ekXAwJh0cz8umenxJkkJ/FQrUqEQgqFo80frXwnV7g1Xd6nNU
xlYePk4v13lZAf4NfJ4g2K7U6HLdwTVALbvoOe7SbgYcY30VR35CISsrdsFFL1KPpHCCt8rYkHKV
E7UNSUSQ7xdP8ijdR1cVy4wdvjvcK0eVBU6tgtSVOPeVoJxDIOOLJx3U63Rx5AbCMvzvuQ6tYc9X
FpOowHPasVb5NgzIbXaHDU5SEB5+fWXVyZrtl4xXQsEDBhGGE2CDtuW9cJeQRB7AhEW3i2lN1PQK
mlesDWdDNCPAIWSkzJ+8SgCzsRmdTWk6BfxxAzliGjHnDHdTQjPylNz+KXjg5BUGEtTg6AzohcH7
QGVV8rZFr/YzB7awldhmXW42NULpAOSsl6kf27eJkBEhYVnR6EVBx+qsC01bcul2eWf9heaNeY0I
lLCDIWtPDW1LAsIHVbhkwqmjOgBn1ERzzRDUke5vHYu5TYazxmlkb3KjDV7844z7GfXGSbgpVWaR
JD32R7at+zQxt3rv0IESoGW+xa5jn3n+/B/p1CVDGMJ/fPNkG+W8Pl/B36OBFyNUMkZ1LPt3cKUg
TG3TnN08Ts+AFnRvBgfBcfmYypWDtOLMLXOWS1ncuIDbX/IDCLa4EEHdiioKFKSXUxauh2sMikqd
Yh+q6EFcaQLZTu6uZ+0hEeS+PhDydS3aqwQBobw11WVXvUJ8o1zE1+IsZ2XjdBkFpK/Ijw5wtGuh
y3FZDYsUZU/dou8hgWIicccpyxlkDja/14RvDeKZGREYzR83gN9pgrt6sVpbf4VBuq7KDlW+omUG
an/M/dv5wblWgkvcx6ebw+Vs7AGdy0dNgRMjdmceo+TmfgG3r9G8yx/y9QVGr3G13jn+99tOjYOh
5J0LLiXhUrWxXVgxSv8aCqUAYH3P5y9spahbcdD9+6g82oDSxeTGzx6ph4/hJsoyvBGV644qqvBR
hgHRUWsh/iqf8w+Hcj/80WIqAcwnu60QynkGLJ8ga+oZGjDv+F+fVn22PVMVJzNyTPdp7+VhfvIS
ns5+8vyJQUr//Z6G6Qks4ZKaKxQKfMlRc1GXl3YDZ7sWvJ4njf+27wlrmgeUpPN1Dm4q2/ZtCuCY
Gd0SdrDDpE4hP9FRYMgWwoadakHb6JORxR6veln/csiHX8VhJTUsIvcoCUBvbBuc4ODgedN4nBpb
E/uVizaeDXnPfVX9gmoZ+bQENRvLyMdOgSgIGwXhoMP6gfhcjxGGCWJRKuDC2yMyJdhqhOQqdGzq
EM/smatEdtGcnxOS4rvD3XT42448pzDGDqoeoShxPu9RO8inQOt7Dpfr+++D6WZNHQocp9gKwdoR
MG3DhJAQYDHsogob2/UxqF6seBjaEoV90sXNHSAgVgNRUxFJF0xqv4FXVl1jhNxuPkVyeyfnZkq4
Eq/24KKh+dvjo21vE/14qYmbo55ZhHvtFHmpoh5Bfs88B3v75St6qQbE/At6siaAKCNia6AvqBYi
z2iwtk9XYBE1XEE9Q7uzuV1p46EVg69eI/+2EVAXam/9tVugwB21yhyn8+I7R0X0YGzTxjN5ZH7w
qxtdjrSE1afvTIC5tDNI5J1NaX7pvr2Vwgj66aBKz2cTpf6jy1n+Lb/IE0OVTkRIxlZ1jI0bPZlS
n46QhDFwwMkP9el2z8O1YuzDD6H7HnAqMekSaobYx5uS0KzDrKmQQbKGnVNrb3V80wNH+Jc0+OO7
afjFppZ50c5PAkm/aCoSfb0tWqRhzvlSoZeI+SlrzOMA791vQdiZikEAwwWi0L5v61jLTK92CVww
PSaXAM2xGysTRAJVY/2tBAGOb+8oHgfrhqVRZ9j0RKi1dCGmmSrPLVMKCaQaR42XIYn7i/SaAVaf
FdBEkp/UHbTxhoPwzFvcex1WSabZgr51eD+avBrFLNUMPOPAwaCENqwKc31Q3c2qtJS8+wxFvmrl
4xeC84MONvZwrwY9cm4N4UsTtMPCP9gYBlonYrY+a8Nsl/AqfVSXQXXC/Ztg09exnPj8UzR0IMpb
UFOyQ5gxME/utZ749TPVPuAB1PUM8W5/nV8rHvwg0Br4VhaZfRuWChBPqMk9jDIBDxDaFxE/14tu
NjVOm0ML9fNA8qDeuIrgoEXkXOfODJ9WfzKkH4y+du2sCGjzI7Ctxc1UjtJ5icWzS19lYgggEpRf
WvXgNz6y0p7dPW4eCkB1B+I4Rf/V2jWMDSMwXeDe5LWtMStit9CyKKecKusLgCeQxiBij1V4GGLv
2ZaZR51K/dBdOoQfTttQWhBAY25I0Qp+lp5dyUvMWagFMh7FBsDdt2hvw/WimXt0eQ54tJ7XVhWe
1BwuEUUoPcl6moNAaocjJyP7SmmDrdTTQAGEWKBG4S9tQ1imTjuMjSeF4H2+L6rH8mx90tkKSimM
sg8Nq/We2AeB0zO9y7yK4rFHQiQTzT08Y45qAiqz4Fo1eESS6Uj+unWwcb74dSc/GqHADzPQl4Bl
QLU/VMpxxB5cOAn4haeb/uj9dEqdoZrkGVAgguUM0lO5wNre6unrR2lERWJ80FynS15BuLxYIxd7
kcJC8IsRyd0ZoSvMo+1JmbwI8YTsve7d578+L65uFHUINGAT4FRyJqgIvE7ZHzQ4hHBrvBp/Q7xR
naY27lMHGvXqrpnYYAZP+seqFolKyAp2EIXaA6USz1aAhE0xJZL2MedF1CEjhVx6LmNmCqcWgrvZ
JHKek04lj5KewnYneb+W891UkplHZW75Kl266kxowOfskALrPcNTnl0j1fpgELCzRnTztFmC9ZGT
tdcNhszXBlbIL1UJoNAmvQX3yiE2Sics09mtvcX0BOTWVcO+QhQhrVlKJAJS8tswPNUsEyzM22ek
fGbUYuuzDrLjVhh4r5Rap3ETydQxc8XoUS+KwGufUuTn5pZDrtLJScw+eLHdU5FHFcvHEUZUWVd1
O+1LphYktXY02sVY2e6gae6G8G/fCrOL7y7Xa0QC9jwTCz+H7UUCcTiUg0hqmq7iQ5CqIKuqsPBM
fdFrDYGglIDW65y0czmAnVmIZjlVuP7JlvYTGvkpAgReYI1S0vL2F+AW4gb/HAuJTkJ6vFtlfm0u
v0ccTd2g7f6fR9DB2Fe3OTOYm0of1/lI1/QrzMmkIElGAOBc7XgpuKhug22giRzJCVygZEmJOt0Z
6ezIytSj1ammdOknTgzz6H53/aZRQBJAXs631AJszA2lJzRAk4WrSCrJaQJkAIv4+HD3nIgvSDtI
28kBbZoKQlHQ7w3aSskRsdczaYY1bGLcyxCaT9O2pfVMdpchbRm1F37JVXsRpCwRpJg7S1Hy53LX
kuz+wEk2Z7Gh2o+6r6i2bz03BxDHok996Y9c3Z1PkmKhUQTcbb9Pc+qKt4by2mx5/6LSbPOCg0c/
dYovnDbZqOm60dE4ZaaPJxxQf4qCRHhj0Qzp1hOzIz1kMEicsk0AhpE5UCEztd/L3Vk9/n39W8AZ
2WZbrBfiV88RyJR6iQqIj/UqnI3cUZ7B20CW9BFiKSIve0mOulGDC2rqsuDfGCOff6Oc3/U2dits
5TVelWcoz4PY7mydZNlN2xe/j8aqp7zEB6K1e++A4MkxGoio3F5UIXfaOXCYKyavuSQ7SYGRIptI
TzJy85JGxUhHCzOTwkii7W9GQwmg2ZlHCQ9JT8uG6wbafvl5FNqAzqmhpZjGE5PKk8C5CNljfb4D
9RkY3weXppt+wX1WfGRn2OBcC+9lsphslru8Nyg5I6hzTir+UPrf6ryQ4hckj3CyyRgBSA+ybpFv
lm+4gJx/ngpeKZZBuxyavHpAx4Q8IbrLHLo4ojuPtJBmeFvS1EvZpFiIDMFwZvslCbpjWuW6jyBX
vEoCmWi/86N7nEONXHGWvZ2RkuaLhyh0qmi5KAfSeqcKWmDS50S6zTNU25+gyaq/rPxznjMbfF4s
jPkiDGgrr68953cLW86LRpMefXivfKx5UaelUB9uLQIPyeJm5x+jaIf1EOJ6ja9iRWz5VLdhFXw5
sVumC1VU+wwX2O+QQcPwBCGhpJhEsY4K91h9clJaaKthi2QC+J4HALUh2PFVoIam6fm7dwpoYRJC
OJHCDdsZmmw1ONxQpSCgcBoRVhrihaqszDm1pfF4LyQhoqsDC2IICeZRsGwjNgJFQzjobZn2Dk3Q
CfuzLxn6g0l+glIdFMeQJbYX/P3ZJigic3V+P5vHpPV9E3gvs5M8+cOs70rwyZCqvUfFqANTggVs
nUSFlCkzDuzJqDFlGFnvnIta9F0s9EQ4f0wyrTKqfOQIB4LXUNdTg1hx4AOetFinKBpk3PCFNqMw
1CzcXI40zOACkA99E7WnJX1Rk6EkJ1qzGOowy1d4Cb6uiiTYWX7wFbB2fOrojjaqVKeT/EAkC/vY
l6iu7hQO72PaCJBC31ftslM+FMGUsXqCNt7J5FN5c5z1W+jKYJbW8X6e2ymJHbMKJ2i/xrS8O62a
FUKb7zYhGONkG/fMvnDasyQ/uyViKCoiVpR9eMl5ttXvpCpi1r6uVrH2oUzT+gRsx5TLIKG51s2T
63aEh6krD5ruDIe2/za1iyDq+w4TuXAPLPcGKq0/kAceP5y4oB2YrCEO+bwIee4aNMoPkEMNbi7/
VquEAfrWpG7ZcSGEpW3RNZsp/Q+eWstnSLGsQ/qos2kzDdQFkzZoSdWhn80leRUohTY9EcKu7ASs
/8M0p/CeyIe1/HiImtA7YrbKnFSRqa5G1QsRw4VFFAOWXYtk6lK0NUdcDKhuPEeBT7U//ICwT/X3
3uH/ynAOEbCbZPOT/lsYRCEtY4wbQtguMCFdyhtlwEJ2WvQCYHwPCG9j/9Hcd0BJ7w6mLZbdMQEu
0avIgVswecMeo0Tce64es2Z9oYVHjb/9A8BAGkU6ENgF1xtvPK+k1xSOvT1lp6TFHmpBMoS4fQOh
nSHjCaoV1h960Lad1EHAwRriq07hKPbltPpufkLU4mN4DJTplb+0SuZhEmq38PWqZEkmsJRZi2/q
lAnLz2RAwaSXgzi3+aqUV34JDo2ZFZaJDzw1gVptx1n6pNfC9wEF4XYkmMVqYThU6/bX1Rgr24ap
R1rymylw4JgMv7GGnBfijxYw4DlEDaSLE5TpQlcxFoHMiIdYlmFR+KyoZNrlMLhG9jge6c0XT2q/
7lzVQxi6hdvSgms1KPtuxQuk3zV/SKcYUtNcOiva/uhT3N8j7tWzRoFFm5CV2hXQDxKz/52RvpmP
xORQzsaNjoU6njduTZ7V3PuzlbglKT+T7oF99az1Xwjjt8siwt9mO95KIZEFDtxXdik91SE8Szb0
5Yut8zuwuf4fdEzuwGTJarURmhy/8JoFkrGk/K1fpWmhSYHCrHTMdDgxJqStfXau5pnTY9bbW0C+
N6m9F4nf8JxRn04J8WiSZm1DqsoN1zQ1tVgXdWtvGimDCbdFUfu5TTAvs0xsB5NSojojxNXguy90
amWr3dAwwawaw99kpIo1rI3zQo9jMPpbzj0jxShUccstVv/kgX6B8plAbUDGQFRxftWKrDDtnVZJ
FAqqZmSAbDPB8dW069M6lN3oFuUF9pozElvAlWDesLGo8iyGw6OMFgW50BUvcEbnzEGoULhN8TcM
dLCJTLcMCJjoR5wuQoxOYlYX9slVSyIiD+fSXi4QFH0D9p1ileg8xqTzNQQl0muDRqM0Xe0Whkej
ZEdDOrJchnARD2PcImX13EP+0tPRiK3Dgf46Kv/cVcOxFJmYZOc0djJFloTngyH+Y7ePrENx2dak
kzQK+iIubY6oWJE9yo2clWYk/h6WknDdOdVxPIJ27Q9BeG9hK96WHhHkpF4LO+U6kPfW1x7HewyZ
B5cywwGCyekvlfLJ/d/o+PrOKeIDEtWNiUPHIKBLyuUtZIlqQuPEFwHiQEdrErQNGAVorT0YzNy+
18RbyR4U/prH/EYjlbxHiEGDzAF+MLlQyB0/yIWvKYtXdMRx1Z0C6UwnU8qPzTYeyxJcxoRwcpvl
7Kn60vnaLyhqwF8GCumxRuZFSwMEuqwzPweJSTfq7ppdMW073QIWmmBbfE7q9Sk3wh66i4ZDCqq7
r9RA1XEwkmcugSJVAbX4aGSJG/FIYLEPz7al47xlUDyGsLAjE7QJcx72nzZiTfN0/+H6uvQ8iZiv
YzYDHvO3j5HIVpYQVjKF80mLTZIk1+ax9X6nj9Xp2sE1Scgdi6VNaVQ7BW75T3sE8cm/MOQkCuOy
VhsuXlmgOjqmMYxep+VoDwscK2jgNUoRB27oqg78Ixtn+PKIlDKHqOKL9tFjQ8OOQEG+o2EZtZmA
ijbqZWmrnRJBdaHEMVXvpO9BGG24O8nSB8wSUomW0DXh9HCrB311ue8fM0Oj/UnbbYS6Wsa2hu8Y
1io9eUxsT6TKlIW4j8Y/cptZsPECnkE6LpESaaHT16/c2K2k828/YLfbyKD7gTA6xgb9rtSABGRr
jpje/MIMsTpyTeK0dgrLSosEdyXk+fmySTG4qu8QI26rpGiZBK2R4g/YZJf1ztp7cuq/oroe/OjR
YCdc5bCT+8kx7IhwRHOWaN8c5xBJvV1pNlxuT8L2k6hDu8WWb5fyy5OXziOzaOBSFlY/CoXPtzCA
qKTE/nbpUQsOcpDo2gih14f8oZjfodFx9WvQRfxCokkjeUH33/ZQw4L44EQhEgTVraCqTNboAKGi
Faowac1PfVS2A8+1TptnTgUvhb6fsTr0ZFexMvW68vkLX5DzzvrwOirUmYyE8770MpsUYR3/+CDE
MzWuN/5XKtR6LK0x+4AzV3mtCWz32y+8F06QinXNCj8MU2q0/gs0cA3x9ca6+IV7PQHo8tHiNszw
hOpIO3w6ZJ7Iqtrj5bLm4Y63fhTb6Qdu8r6lPZBB1gwXG+lWnQYw6TCwaoW7fBoNRdM+FuNq2uXs
t1K8H9l3/X9iCiSV4Fx3bulsxoJVK4VWh3Vacn2GTcJ11GZureG4MIFaUKS94yP4xXxxds7qf0qX
k8iQTaaRV0ce1d+F5lBu/D42vjcf8/w31k0hT8J4NOlueDtg+SBcaE1SXZ7OxV0BShTJIuuHjRVz
AhBNZ8SYqcpY0BLT3kNYEp862n4Qakpbyjzy5XY6YDGyJCwls0UlIkpdMqQimbpFKezU/TWzZ+gQ
UaN6Eh0ZGNbZcEV36KqxBwpjkXlnuHja0rS0yHwfRt78QqAtfN5obDbVN0PQXO7v+d1RYPQWkJAN
j35lZ6hPz8zYK/URmYRgdJn64qP0lkzo5tMT4ZYoYXq8aSt/yq6WAbYtYqbweb77kEivI2lZVT0/
TS23wWSpqPSJ5bc1fu7tlFp8MTQT/jTnJJKrxV2zm9PKU0zzu/jL+ry2Au4XXc0VfnjWJEwgOKj9
76O2+hWfMXz9ud6RPBRU2qWKBlsCWMCiOKfIzArybUiZJlJ3khp+U8HqOzvxjflbA3KJWLKkaNG3
weBw9gkyEzlOxfHXlm5tYq8uu+S78+3jV7m+Z2FUVYNKOjZGtqHGlRZoBsPzr5IbBP/00BdWRMQK
NoSo2E2Ty6RI/SSdhKkVmemOOZcyUJ1adWrxyHVrcikgD3aoXfVWLbS3E0jy2fl6ia0wrY+gpFwK
sMDSnHZxMu83k3+R/MWmA+5+nakWe+TvSUXiy0jl28vOyKASdbPyad60eW5BUMugrEVzwM8m0zuv
Af3gIwcb7Hkcch/GJilF6xcvPtM9Sisv+LgB68bq8Ri9cERdoIVcTYkfwFpeXhlOLgQgL9FZ3tjp
+FthLvI075UTXpOvCXsNigML8tGRQE9dkuAbx2OTT363hIWU0W2bM8bfzQVx/tZ2jGfaBjXUn0S4
7vaXH0nxpwZCXYxXOyGDtk6PHpirX27qOEM0v+H/7ro6iIhAiVLrUhawFmv4N7rr1sraECfDIH25
9Y6iNUS4FgSGMb8bujwxcyWgmdOVZMwhZBU//6DnEzQh/Id1pDDgIppQ4lIitstECWHY9C7mOJLi
fOF8fWhzAVbCSMgVwiizVgMsVbt83cLk8Qa/9CT+d7+DZOS/rrEsehc4TONVwv8wpsUaUVDicfXH
Al+uyTCwVmp1v3fHYzZ2fh2UADX7FKUNff50fbZTPwnTz3aqV0b8NSsUL34nEkeqzzawdfuGdT//
kLkDqeOGwvh/OFNjgk5VGC57YpXDeku/fFKhcNIweQFVGpepNd5SSx21er7z4V6oVrYGxGXSXNtX
4G61J1L57uUQXLL0WusjM1dLHEP0E1JCW7f2AA0GGY5XQN/sEwfbl4IcwijG12bSP6X0THKNu5tn
8n1CGlNcFviaIe5092ghq7wBctRTc9dtn21gV4ZdbFy6ZXDkrJ/fDq5g5gUPCyaS3lKNFpo6B/dX
vzGRKP9Bg0oDiSWdzAgsSyVVLYqqj7HnEBzmA6PC/5gOnh+u2Sjk+PsAOkG9I5oqDw1zkAOavvxp
d5kPfSvv1MSCTEs29mACz6gYqd4+6EappPufz3VcXRa62YcnvSG90x9E/k7TLneCBQnoLPKhTG4J
GajieKxYyODCuVkUEuSOv9pQoYLxiNbm4+jIH1pV05PhcTz0X/UaA7oYrm7Gycc++A8aY/ixaadr
Ij+n195AsmpQ3VusdAinhSNbbVJpOn6pnaNifRcYKLkyjmr8TVHTzk34M1joELz9yM/6wBI/5aUZ
gnTXkfyZePhMvF2XcZTm1BkfMl4KRT3FYQRb01lBhD8wf2r0r6W5wm4m4gXdr5hCBaIS9dSUkaUg
2g6HOuFoG36DB0nEpHCXYPYaR/Oa9EEZxP33vkMw1ekxT9t1GW7J/l97OILzhnctRAu6CIwWVVAt
LvbNTtUhHso/lWQO3Ry/olkJvsOMOuIuQD+aZh3D04Hv98R7lH+TPdjzCGFGMPFmwfH7VqhZscI5
NEAeUDLmL4J7ZPa7QY8CqGVJdSybOyueQiKbw4liDF5f66KYJjRK1uG3Dlq0XeIL9qwuRggLnKyj
EHysFl3bSp0j0gz0eeVeEgy51yqzQ1rBKxPUV5ivA4PBb7dGYkx/+JfGGqDM4XS1//3kV9H5N/F9
2rTzZ6nds/5O9Saw5tjxGRNsb2QYOxcpV1nsMM3Pv1Cx4PX4AHIhPdDJ8MCrLywaWvvmic+MB/Me
qYER7nxnQUed5zeLLYo9yqzSYQPcxZJPSCakG/x9pyRat1RLR92e9n74ZQG9exfnpx+ZhWbExN8S
KCg5AEW+lv/aKq57QaDs3uOCPdFm3d9AfMzzLr+dzS+G3mfFMPbqfMGdbpEWOVPb5nd8qNvhNhI/
jRnjEakpVHqMTbrGRXQMsAd2wMxYnnzDWU7qIONsuPLp7PPe04GeObZOCwzHgRRrfVmyw99fYtkn
sOJsrdWJF5GLho67xQkm4lvIrsnpaBkgo5hLAn0huQLKihxdYWF+0Qm4xRsxQ3Xuz/jlPmTIhDpX
Z0GKZd0kgaHvHCorrPDfU+vljE4AD8k/poTeCsMB9MWsvRIND0+0drJDRBqGXwFanfK40KUcd7UH
dhC0346f92magGa4eNWFK49a+QiW31ieVTT4gDGeqoScxUVhhKNTpHdA1ncrtaB3T/05VY9dRLwp
3ZSmTh7ZXGFyFnVeJwsDSo8G7E8GpcQoL+rcQiC8Ee4FH49k5LP95FE2hR+Sa7qCdlqaIkACT6Bd
n1GZf+0GNPMtxWDDjFt75A4dcQNhQ1FYG4h6pCTbubEvBMAAIQ2IUyMs82E2aGTS/puVWFwh1DcD
gb2Bel309niE+oMd4mzqxJVElFVR0iw725gyAIUYGPweFU0pjpAH8NZdRtxjLgXgXMGl6ZGCZpSC
BwFZ3gIZw8QmPSXe1RD5Qi6YLJubSHIOCDJI4TjOHka6SAG4UzHRL/aYJIqAsE9vKZxON9NpoFmc
KGDG8lfLeHFhK0crF7SNoPl9FB3sI0+sZGOaClZi0zDQkOgMS4SBWml86wpDYGv//YKBb8IffedZ
n84CvkCbQgOtqOLARFFBIMSSpvhZSraBWXCj93qcQ9C5nQv+V+EgAAib+b0/TRxaH8mwu+ht/WGJ
Fy2NIP8vYmDx9ymJ+4E/CiibbWP8BaeDqACWLoo6ZaRBwP/15uFp8msRQbZHA4HOW8q+Fo+sn1vZ
/oGExEzCm+GoozN3/bZOWuWEkgtQYZnE5SIgRxlvstNyhqOp6Yl+ODyY/XAXeBIMT4GYLxqogIlp
99087iCnUZ30e7+QQiN5/wTr4YhyB0qBhMiSSmfdFr8oFv9cFA0PKzLKpjo41ILsrJqUOMfO7Zkz
QvstjkdBBrB1REt1DHvgMusOtuYpPmKEdw/AYyuJB42689BC6rrr+6KW/g0qFzO1Q8857OoF9DN3
lHlkI7Cr3SjsVU7LFPIZqVBL+BtW1duxBcCH1+RkDmytunmU3YieKfMl1hh1OF8yDPPKRarU6Tkx
PlKm+opvyrA3f6NG/smJ/TCdHACdlL+BW5ec2UDviBvbQA5Oo7yEB8RRn48fmDZZjDBkFvEye84z
BD5s0J/LE2geN2lBKkOY79tk+cE8ndbwbR9mWPNK8oKuuoP6GT/yd2zLI69A19+F6aqQWTRLYs2m
0rnE9CZisk4AjGbA+cVDyFzpDaKqaS6LiUNmO791YKBv3QNqaF1OGvRg2dCMN2MZOpb+5vqzIZp6
XB3e8pjru61t+i9TYIaFbjc9PSTqycfUjhXk7TzKElVP3MSsCz66P1Dwf3t6OAazhAGHe9bOBeOK
qcK1OyJmJDDmRXl/X7xuDwcxNE4WDLcJthUx2puudWrY1j/X3x5RHGmXGldNdrhf8nVYT3Zy6aL2
bmZcjRUvdO8NUPYyxkldeI8FFZpAckvTiX1cYZQBvPjjBVQA47NXQJFIeyiunGelrd0RshEYAL7M
WO5xN+IuZtlj7ys6eVWxeECHwKpIu5DlElW+fymiwIl+YIO0Lz/LVdrWisMFAhRp/PNFn+xe+ZXj
pH9yKiqP9LC7McZ56YfCBS/b9rnbLgQa9UFauQM/PbQokBkOm1mNb6BGtrlI56zCyI8j2RzJkv1g
9AbxJly2kOF3xswmmIYXBTYOcJoI1vfjquNAOgRMaCFT8sdeHDQ/wV2Vf2rC1Xn3xnivrC2P21nw
oUMBcKDAPRy/A5YGUS3DQheYdokmbkw+Lxoi707sDXtp2TGDJtZWBn8qMYvEorwlhObIJuiSrzyq
VsHCp7HVvzxE5WweZj1T/u30NICIqG8PMCAcNuEA4D3up8NPN9J2wuHPMrFmhVdoxSQoC2c+ERw3
wbf1DSdV+++iO1HpLONmtsojZQAwCqsIWQ7UJRPB+LGn5wgLh0LIpderwjAE2pbNHTnqL0Pc4gdI
3oGnM1iWa5NhqjiRLxgZBVit+c6LBYO6xQdR0KpPdJU3mdFo2SkHtB6m4mZ5CndxtKQKjCzXyNj1
ZIj4KNgucaueA96qbXAaCLejyz4B7wMRToJhINWOlYm3zKKE7JuHe4doLJzD00c1VYQZS/YB7die
oefHa/Rhzv9o7xMpv+NSpZVQQG1Z3S3xJXr5jTcP3y6WZ2B2rpMODBy+L4pMvvMxOiZzEJ7I6Izs
LefMWopmcPYkNbIEMzBw0+mv9oL6VRG1bc+tCZSZyBKT+wJGt4es5dMKVS8HrYQ6HLgj4FeeBZQu
XSKltnI2ZAMaYZCjfJqcJMN9ifU1ufpYN9tneYtdttqPOtNZvPFarnWlO2HjrveOEsNGwZ7YCFbo
z2RaiDdtWO08dFqOeXdu4Ft0ylNyGH1Auj7Hz7Plvxg4FRvTvpoq4FcXI4y8/1csyqLbsmPrHd1T
WlU8XZ6Drb7R09swBayY20fmiGXUMKwlYBqMTmkFkR4JVpk58MUdM6sqOm/OlRj4N23K+UJiR+US
bst3u0Ry6DuUYZi4MN3LvZ16Yc3Q320QCBPn7Zy2/jdG7U4CTrgJAuQ1tJ78p4ZD0BodAn+oHN8H
ei64OolT7DDy7lTeadIjYcoQ+fqDniWtLYRlixZljY0OdnZQW8SyyJsrvDfDbQnYsyD8qMpT2dpQ
BaLEOuoZ7AboIZFsVbR7aC+xn72MJ8aZh0Fy69fLIKJA9rHkjD9qtmiSu10ArJfX36Hki4TuKuZv
60TG9xHkT4EC7Yxcq1ku4ZVjYNIobyCTImEZSNYDWXhWQByRZmWsGTnMKtqM2sees7BtjuR95khz
afF8UmbuvOjXJg9FCrIZT/BEaUUZkb1FilSnvJldII/tDjzzG2M9HupwwgZeccPUYuSkMXdp9ksy
zgYQOlvhlMv0ymM1AN8vKojh0psAM48o0WcyJA7EIYpYyxrdvg0Wkoc8Zssx8NSJv7bdCcoTQqBl
KHF/01ryUX6QryI8WlI0+mW4z/Jpx+lnGEHtoj5AiHZxmsEfIvb9DGmNUfTEKLO5VNglRJj2IK+v
xcOe+fRYJqxYnfMR9/qPpBxJgm58iYH9vs4L+2/jkCKbk9YLuZS+/q54ljVRNxB0ZmrSVR8noyBL
UZz4y3ONayhMjFOV0prYZVGktlB29qHG0c7zGFV0qKzSGJig4YAYMAy69RiyxVLR0K/ghRVP4P6Z
ERgLjlFEYaiUSoy1ywdl/jNIGluZcJtDnl10KIvNtBPHCG+ugMfe/O6HzGRfL9ii/wrZyP8PxbjJ
orsI1k9qUxuTGFRcO23nOwBORWIH98oE3MGGmDgFCN0iPe92oCrpilJxL5fIi2mqfDxX93GPoy6n
wuZz1q7ydyzzdLwoDKXDlwIoX/+rfzKoJNPkf9eRvILYSdt+GA137LXlr/eZqJabB6JTJ6E8dR9+
lEwhs5R5Bia8QNFxwS4SnDYfQFpmnB1TtTePyfn4tBQ1FPDjzuhoNQwL09R1ijSe8sPU6JpdZLaA
sdYXQ6I9kzueSLauSTq+97RnhrqVjZsxEUmRjcFaxqfBd3rZnIy4iWNNeKzPN4UL3Q1fKoQ8xNs3
UL4xSE3EhQa+45VLyvaID0LrDAMdaKz+DYE3PY35TTrwA6sK2mw9sXySNdFADr5m0yZ5uVrA2Jnk
jIgR9Glp7gLTqG1WrsvkQk/mmag/tCZGZQXeBBZI6fUV9IO4If5hg/ZWQkp0M/0uunPyaMyOChAz
uW592+PKSJPXeJvXhYPAIXFe2woQn3eTgDc4rQHyiRmxubz0/vVBH6b/hvPZTV2e4RiTpH7cgthc
N1se27vltyp66wq1pZTexpxJYpOnEXRF9qJc3YzdOGqBAu1rKet1y0EBsyY1fNa+AM7hNhcFQ9Gq
NRaeFWq4d2SKPCNCPYSlZq7FrvQK8ijUwCTV0qolMUxNRg4Xs6EWdKED5z1tChO4i/HjSbpdiomc
8OY9YRi09/nrHR3ZfnproYCNm/n5k82LWiGwLwvx01yo0iOgxoJuY7NU+EuWTRubEOBxwgJkPgY8
OhUh7joue1lwazh/Qnw8XeZ8TDKxbG3MYt1unDxm4uiKCEMe61nX9mlfpBXTPiPOvxMTkqMeOkW/
Q1Vsx7qhnrlnHtwU6oFC3Ajoe+2kDdHcCQR/SAXIcEfpPpIOFUmyZ1x45oHe2A0rpU+1iAxNZBM5
9Y/cPHHca/idHpwohEBapruzEYR9q4G2XI0jgqaqQn/qand+Xh+Fm04gf5L/5pSujtCDCRLhkokC
NO9alNLL7esIUJ1kFWMHhHA1acvAhzl3b9tULwHU/N1KLaZlhSdWwFu7Bmd4UA5fhk6e8FIdsyjm
iXxPzREeUWen5PR2Rpfz4KhKk5Jib5ZxwSsStNb4I0ThhfljYE88D8swFDh7Si7Fv++JmO92Ra0P
6OjC++Vp2KeW2DcHINtCCsTWr8EMa5ZhQFZ3ixGADqBoFd64FqWxp2Gsy9mRbdZTlmAeFmqYoUz2
kQnRpjGPbLzYwY0VJdKP7ovF/o+REbfGdD0X06NA8nmIgNO5Dc3WNj0r1Bi5H0rc5d8QLO+oA80h
hTHoilzaKFcpSTblAC8SaGdd8J++Rq+Ui0AcsqsbVQj2X3M+T9Z0vfK/650wJC97/mEjEwl8waVe
Flu4DfpVfdVr+/eOj1AaWQgxjocQxQpGH9Jx5GqXhPpJ4t0GN2wh+Am3GQZdNeBxzGis/TIrft50
n878sSfnwYZHwJASTe5w7fdnB0IEzerasht/bHGR5x3CVSl5de1g2huq6mXBv4Si40qEIYuMAcca
N8JoeKi3JkF+/SgsbeBxzLdUM1vpPunj+M6DiK47eKLHaPxssejZ19F4HPOBGNQ2XLLxqQBohMkL
fvR45VzvE91ngcDmpIIlpTjdrRRi/Sbsho6QbDTLOGKdgw29/Z2Pagrny1Iq96n9eUBderZPUU2q
n7rpEGk3QLjHTHTED5nujr09IddTrd1C8RTr+NM21xOc8LuR19TVumpWl2LY4KXpiMcwoU0ydXLy
0vdcfzvxeYtL3vYajbQgnadLvFl+S90WaT9XNu71+fXEVtETbOCbmY0W9Ui7Jq9jw29eyjxXGIzo
jYXuVRoxsitWTc5VpFjeIb4bWUckL4e6Ln6CxEbNthflz4Bh6vi7W4D03BQPyu7ZKC2uesCbm4TY
bLXMXeahZdv6bTvYXWHAjPVpBPoqyYcGzAn8ba5UjmShPgGe3npEfscfd+W7JGBzFcKFap+c3fo7
3mA6G13pdgmo1rjTpZxvZVN0ydaXeSRrC5XwnAHgZPKDwjREIGVGvREv9mFHaQm2SOzwTb4KgtKN
ZrdScd4y+JD/p/PaVTf2q7C+mdyf+lU4DhUTlGb5YJL/yKaEgUH3CVWvwLC/6w1uRyajvL4YrV3h
w8L68blA26tETNq4EtcVe3SWvoXfvujaoGHsWLNoyhmifNb7tYf/2lJ+uzkTntbdTayLYkNXi+9Z
nAeglaUZEAyYL4bzcUAGDvzzPi6KMOCHh4jYBvjlvwZGsBfGqF/ONFtxylbK2MttlHChShhzz3zh
Wp3h4I6fUvfNZWhT80ij5Qe3c/VesaDyYpuAMs6xJEaeBAPyVtz/QjKWHrGhZcRpDINjnybrsll5
QZvYdp69EXe8i3AHJAmqstM4C/1zvkN6zki9cRRhnk8vCylp7AtbR5KVBF+oDIy1LSJ/LrjbtFMw
nw54MS3HpD//jSchKhm7xfVAMsQFL0PnMBShilJ+6jAc+yq8Byuj/icSsXMr4Q9oYBdjNkehJfbi
YP/d+LBWCeCxXBf3NNG3VL7qnrnp67YxAHR23rahlM+Opb1x7IX8TGDcIzChV+JvYGp4IZwKc5gt
Atzk0DtHTYnyXSO8alAFbW0KimEUf7l7J4yL6yLVaGH5bhB9Lu43ETOhAHcl8eXX4br9locKpdG3
WLMXaQ1oyxKjPA0M4F3NhZvmZNrU2CE6aDpV+rqUZaM2yzaDSNtxb1eDw6RW/1x3V8AQBy6FVY47
Ej+GzD0Vbr2PzhlWoYJL3+QM41K/zogedMXjs/YXwWVbwIjdcKBmM6BdxEslOLzmUsAm4t8sZNrs
9ajhtLtfDZhzBK6nloCUF6MATIWWGF1RAzfPKBgboKQMQZv7/Zfkbf/wNEybuWRm4IychsDer08L
QWhEynKv/SUVGP9Jmig9sk1Rt4Q4i669gi1P4aqM+uWyfQSLJrILcI0RP6oCfpfGvFOulhG0MVCW
mA2wvTFLiKLp0FITCF+CkEdwNdXMVu0q6cuFQF9pYqq7G8+PWLuVnWyXNw8KXiyoEYpF+poYMain
zyzKbioeB3WxeFbqaqv9S681RGAkI/JdSHpbZhcKdAXfPZNc5lHg5+qS+B8xUcDUAINIBzAoBqkF
Aaozbpr41n92oFjtz5x+KgnONf+nWvNBBT0ku17Co3qmVd1XBND8djYJkZr+PO8AgvaVb5kN8nXm
XqGHVSlT6Snb/wHm/+5mP13ID1y2E/xGcw2mO3ivDJQn8vxhnlVyycTBaEaUaFsiFt0JkWeSaXoC
Q2dSiHl5HNBswL8yh5E04zxlxBmCKPTpHEpRM3QbyMG95PBC6/+5NYtjFmbFICR9wD7fT9GhsgGF
6U+sANVry4l4fj5RNnjjWCYT0kLZjgm/+KPaYVVC8pg0DCGqFeKYXEPgcVjRBHSc+pBjmcHX/rrD
6twP+8BllkbX4JiWUySTsOIQYB0c9wISdZxXpwtChdQXAi4WztQLJLgTXlPm3zJ1Bq7oR9PnYQRI
SAOFLZ0vCVTYLrNXXzjUbk0wExBDyildiqCiBj5jQEXOBmkmo8W8jLr+33nZVST5GOtaywaRrKMZ
dIFEZdqrtxkt83TSGmBOWd67dpYG8h4BoCU36+afVX3DAOoKpRa1Hi+6/L04pkX3QGniPgGnzfmV
BLWN/Dfsvak5aoUdu1r8YUhrkL1uSzdXfwUiooSUJArxFBI0jAqvexyjkHS2rEXfq2/1PSa0559/
G2hiSq7XWEhDEfqsn93Qi6Fr8/S3uoSJ70QQPZ5RGT0PwIBPtjfQPTFR363HvcyWM++TXM6RekrT
11vAIJq5kf1wDLk2oDVgFyHQId0XHcPxf/Aao+UCvdHe8BJgAmWXs46V12xse7XjYHwWwP+pqP9+
NaxPrJT7/UNUXz9YFNtJU3QI6rkL89EQlD7YUsu4Qmtc1u+NYSnnDI1fB1UfcYHRRk8GYyTw1Vyt
TC+N6SHWA6TVojKeAr8DR1Bc0MbB3ywIi0kFYBt17pl3DrDpyLvaI1CC2GdMc38KEHIop+axwNYC
WtiDv1/LWMoW1Lk1w0PV1x6Nw5nZPFKY/A6MjheQfhzeqdIpDtJLNyE9zpO+goMcuA0TxekGPh7a
h+H3yp9L6522LvarXmzl5Qkd5CHCCkiGmakG3bLgwzrSGqapbWSa3x+1Nt2pR8AoBmS6hdGwivu4
DNRZC9B82CJ2IhWSTmPnesHadJKBxlBNpqyKb+RJ5wByOvee1rhtRTJNGh5DJfroShv3hwmXsYd8
Y+sZMPDtbk0JvZifJ4MbUpdWaSvgvePH2vvh/lVjiD2PK7ibuvS+6gUa1BRam/WxpR1Ob3HWy3Db
9a5C4gTJJL/w6kTwfWIbERDkFdwi9ege7Fp6H7kHlEqv3Q9JGfMRFZYHmjaoQhbGY5o+g9eoWX3K
d0eWI+dJxbSMVdMrk8zrDE/Z5xjLr9jAAdxQEDmHY6H93ckKf/fcSjD07a7zc1Wr4xum6eYoJsU+
9gdySy+eJ3a0b8v5aZpZCPdS3erZlFR6vOjvAwqX4QLzhqf6qZHUTDfjyWsO12h3MFJV3Opof0EL
8ZhS+ZZ1ugOQzyDg8EwS1eEP1tOd4r2l3A2KsqoGFBuYX1JVUXxnkIhlV4yflb919FPfwZFc9VEz
gT1p7CQEDKoXKn1g3WNukaJ03UvTYxRM+OVv/dw022+uh8ANAOQw+POBVsDJT1GrdgnPBd8VqHQf
T+E4hIWjU5cXDkZgmOAgSCRUiwlh6+NBYmlFsRg2TxuL3QXxteXd5gM+qJefO/fdz0K+ZeWoTAxl
PGPlE/XOmcd20OloOK/45ppKxyUcCo5dorcm1UApvxkclQhU2sm1xXHlsXHvP2bFQ3xUIEAVLt8m
obHMKfSPi84X5hJfI96os4WHnhajTUZmWZgRjQDDQPOmEFg8FIipjqTbnvVWKFs4UROcrJNpkeoE
953XdvS/tT0X0mtauXArQbNtFC5gWE6Pe8s4N2oGMm7dPPS9pZ/eM+YugjK7iQ8+HSoXT/VjsLZp
gpmopNVy8VpbDZewVe9iPUbr6gpa0fubNqPo+jOsm71g6EvLHnJxBihXjyPNgVKaUAklgHZ4Y1oL
oxKz9OGUlE1Y9CkgQL6LQtUz7qbOzxRNVJsv2TmqbeEslHAmC2IgwbZGwR/h4LPY2OZG9wZ3YiS5
1Ey8HAVK5zbCwzRx5SDAetXjoms6b44biDRRHsTNPHOOnQ120HQuTSHxmkWW/y2VFxIDl+MjLKYU
BiF8vW+greCP/9hcj6Mwxsgpl3nxxpfAgJSe5PHBXG7n6VN6pyDtRdx8HOSZLw8UIPQU0b8GPuKG
tx9etglCpmHNgEU8vUUild7Y6YcVW5thgRIFHn8JBNEDz3vejvE+Owh9+yTQe4x2iOW/lvPMeyt1
Fr1YzbecVLCwwdonliLm1pCL0fB42DqN5P9p9aD3uOdov0FSfhmjO4QvDZot0HxqELld6Mw4UqmY
WCodVCwN2XeQ5rVetFef+P2hgNvlpcQpDgWEsSaTLb3igRZMnCCTc8DVIW1rnMI2wINPcu+3gvf9
4ynu/JLOSy1c8HrgZnnV3WZLWJ6dJVN2+EeL/eJSIAmX5HWAUchTiht9qatN6MsGeqNXKxhjTyGn
t1MLTFYKQItJQ+xsif1EJPRYsjEHkOy1R/ylTimgWSEmix1i6vTuEoYURsuDweXFM3qeG4yeO+fh
xD6UB+/1Gk20//sUONVNO+fLW8+p+pc8R95j3TwXesRm4Q9s57ErsIwZobYqlbR1IUVo7Y/cz6V9
fb4BzwAIlf1uWFYIdX4JI5mI/ZBmHe+Ow6druSdn6uN+x8rvIiDG3K7c5+4dz2uArpFg2Az5ioym
go7QHbGh1nNab27mQsVj1BLTtpgxcW22DpHHOZsBLgwgr+BuC+Hm24h7Qe6jPt3q9AR3v42INIPt
cP+rolaGo8gfsdB7esIvhjwP4iAUmVxX0EuQooho/ylahCm8CSeOgg+WMptZNFGyLhmCIPmA7RWs
iE1Q6XJ0H2DAoDl0ATaOo8ybZxgDBGFmvW6T4X0pfzuSaAWtAGMp9+GWyBcbw7uFLzAN9VsCbyIB
pwlINE9Qo5MnJ9JS0mLQsn1FZWFhI40u/QrPulKlwR3vuqZomM+jH9vix/D0xgnDZo+uSD5/aRL1
B5ggMgHu4gR6QM0E47Imw2lFQ+iMLZNV4XQWjxkWwukVeEtmtSBqAUIFAJRbQPg8vQpEa1m+a1GQ
oRnirYlT5dZgsnFLHyELxR+eSZ7HkucDzninQOdFYCotudOkOYaz8uRqPYYhIvAPKAyKGpv72mQx
K7XlMMge1oVq+tPVys3FT/zoYEzG+6hZAKESh+54DSRH6PjEzmHuRyUrZBXAaBDLyKM1OEfeTuZx
2DcAb2oq8YYU9YdjxH7+lRW/kXv6z4ScKUhXzDXIVAjqAZAVOBSS/DUMNsH6bCavNVM2DOYMqc5X
CFNAjr5KHHUSP+sZ7lOuviMsSyP8EiE50zFXqOJfM8/TBhdUsGs42P5t74Eg06v1qe3kmafjTGza
5TF646Rhp30zuvCp0Q04Mrk4kZDe/K2fyPh/CD2oL7VOIyei7tZibcsUQIW+2BiWtk9gv7e5tgsf
WlMGXoXrpudjzHwYmcTPIKVwlYhBsiM+fB5FKPdaPqiKK7J49+9benvFs/DuwgQD8ugKSt3gDAt6
GyshQ2q3T9bWvls5Zzi1sB+1Q6/NUI+pflCYmkwly0ZGMXH3uux81HoZFPieoHlL8fxua0T2WG9i
gkpltoyY3evUeaIuOcHCZ+ijRG4jfnuKn6TTgQtmDfkP7VS8UgCwf23zksSIevFGsWuhXhb/udWl
S7akU3dp3eE9LYjoD5IuZd0yz7zmZX9g3RisN/JhNA7bOLb0d4KTOPKXW8eT15L48czeFKx9Nsnl
mV0er/o4ABE0smXsIpZVPwWdc7GkyS+oGWqkyadL6ljNB21Q1pkrxhUNKjYxlstw5KZVVH+wAi0R
Dc6SqSF2U0sMw4opihRcZtYUaVqnLdL1oEyAy+9mjAEDwTS9+4qXm2bPU9+C7LuM0ZQj19YWF/6c
TNd5f1hGKXTHhn39E9O0Re3hv1TgLp/F4ER1uMLsQ13Pf+mbu3+UNrP2K81OGDHavn2Olfg32sID
2mmY43voyUVFLoVd+v06JtccPq+Utn4qocql5+MM0BrWYm2dvnoDeTnNMA1m7iecVKMr1GSqxeEn
QrXnODlmrWpsd8+oXnWyRwgjX2r3DAS+4VpYJrI1tMwbMay5JtvmSbpoU3SwYRvSGRUqnnNqHiOn
iQO0cv/GunqROFxiYoQA1Mlg1/4FRnXGPd18JkmOCJApnIO0SaLUmOlQQbUBn9PKgJCKdudXlsBc
/1wjIlWcVGk0CzKAVI5iqpdce0K3DaSOd/SjUs0HMc1PGPT0BBmleBbfH9kNqZZda+DxHQGQsr6U
BeVtNuhHPCQLVOnTXzQLeiK7bMkDrMf08YI5DCwP1RR+M9N8Ho+DaTJrpRrVcEc5weOvsGzqIF9W
jwOvM55QtOUgK8x0S7ZsAH9gqcZKVoWmqpj9zys0OGQHXyXoPahISiTlj684U+KYY8vDxmiFLXwv
aksKHEkhm/gxTWd7FuIn8RhMa/qAy9epXP7YA+6c5JcNtAs9ygVEU2XvhIqCDuwelzTibatAz4WV
FDklS60W+BTT/yl7/MZ+7bWTEOzaokOsyIUJsNc58u6XxD3Hk8OeEe+NkNGGBUGehU3hATSZ+GqG
aap6uEEa97eQ9lpYqynGjwLalvCgft96Vg+WU8VR7JOqRVhFuWnP7Zsrp37OXG/nl2+LsYrVrSK1
yKexwy8kc8JWZbuHojS4IA+IO6ly1z6JfdDPAGntMWi8Xpk/yr+GCLKhsiCY4tVb1/avfbX6ZeOd
wgA/NAr/NNxUvNKJBeqpUcB/nytO94g4fK0jQPziZw2upFvtysVeKlAGeX0eWrEP/n9M8y3cZ++e
x7v6ZR9UC34QRVeV5PBt4CIvByCUtmZP7wIr4OIk2drjM9ZgEbWB7zd5JrQIfdl3zAkKmkeHKX4d
TvZJ+No/Z4pnccMXVrzfM2pAipc4K3kSapyP0oyKcvVOo/0foEH7oYpcQKfc8pWC7ZScVgA/BKF4
QlFMfq/XoUyqN/IBdLbQjgoLO51eG4By1DkpKe6qNUdyi+mH0BplsDc2pKeSP8A8VsszWGD33mdG
2hSWsXCJf/NcI2b4cvN4CzGmt1AW8veM74eDJtY0UMq7zQVYZq7YeXaFEMtvO+zmALohLX6KHBlc
ywz+K/CWShcgrQVpz/ZQk1CS1bGED14GJKfdbNF4fK0YpiN3hFMMfPz+u5Bt0NBRR/NyIK3+c7bp
Lp9dssBq5qONFI+bw1RDyg0mAykFgLUM0qOChXVtAh5s4MR0/N6M9rViGyuNUDQPO95oG3NCyHO1
V6E3PSrWPP5qpWFmDTEPG1UY68Ij0WL0+iTCsph5EIPZyr3NV9XXahEX97am6njEbahDZ2hWico/
CfBOG7DOuaU/qj9xJIYCB7b6hi5nt0a2LF0uDwo+iksIYvfNauodvekUmDXjfTIJeXF9S2RpAd/A
MNXhu9T3Ls4o4gl9L0obC+49P21DO9zfLaho/NHmamAhJyR1L2xLHaHRVwrtIxP/jBrowD012O2W
oDRoYnMgBtmCYUgwcgctFwHa/KkFr93iDb3nVCF/lAe0V9BYeA7P7uBxG05kK0TcybfGKXiwdS7h
robQDhG1La6QzOSc0+R3vCFT+t/LosOjL9iVZ378ixOfN2kbyfKb7LylLQSxKNsghRTfYE0gQ6xP
zSRdZFOHYI3BWOJ5t+8BMFWgIOl0WDBecSxFfCsUIMaoEdrI88H9WWrA6t4Eci/b5FFpW9l7bqO5
ZzFvomwL1YFlnCucohO5iT7OY2poleHf1l9k1FCl08cjTldMGbfTgG5vzX37STXS4jKuFbbXTsr/
OB9EEnBxOtN1s/vM3VebiQjD00FwBTRVFnDYOBm18VCmLHFV4A8GbXjRHYima2E7t4K2d9l0BIuo
k2r+XNGDUYYRFWzlYLCarMFxKls5SZugSSSpUBW3h2wt4W8zSK6FHmnnisH8Z7R+pyRTC2SRifAX
1JqL62KAdrf03aUjPxBJCY7i9sT4u7IZ99HpmPNMyrZJNzWFjL6fDA6UZYFRKrnTMJUOsBixqtJz
5Ov+VsDAuJ95eldENpmAkac5UCy9AjA0y22MBdbXDQ3NNKk9tB+K+u/XK8+nNSKqqKCvzAWcyiSv
orhXVl4SeLxR71eIwtCdRe6XmpyxY23fB/zgD7Gbac1LvzE4bQt9d5Ak9iUAahsaILrwk2X+pvsS
aYGRVRKWWgfOZX2RTdbP8vSZXj9Pk7dbmbNID6sT2cZ7CDq4GMNSJ0fcUDVnprzlFtdVqtSf+3A7
9W2qIcFL8ZQglH5B1sQaFtqdBFrnVG+G34G9ddc0z9kxsVbtkWAW8SjnVu9ydyjSoIfSUdCVtLmk
s2qgA3kdarnqLRRGPSaOzfUcxpwjYQ72n8Hc+jBG3z3exTTVgBWuUm0Ma/k/r/Jn7McNyUfdOhTT
RhGOa9mmlGp5hvxXly/m6WRo6E+JvhiqQLXKSHXUELBx8Y9xayDxSav1PP89t1eRXYWzLp5hRG8x
qcxTmpFHGG/ytc9GGXf8XQOGhp3aFu+qIJ4MZFIQP0tmLxp2AsyuhctLZOX1p5hUV6Tm5j/dFX66
wUsnU6siMeRNx5ThbF2HNyK2btbqDb03rD6joX4KTtuT1EOGVa/iGjfOmEdeOgLKUTOdsXRPdMeb
CDOp+1oswBordgiGK7/owerzIoH0m00r7cXqTHAoxo+Bt+D3N6ubUrmk9xm4PCudpLJDBX1d54sy
zvi0Jra+nlQA4T7PSmJAFBAzhSissXLQDvgF4KPXg6rVqv0xo6nc7LT67E2QQYB3mBHV2rqiZ3ll
hElG8RW3yB3JTHVtFOm9IPaK17WGxIRUe9VuAsxknZbCtrs9CnTMvNYNgL38mdDUAPBwZsusTHFq
0f09ZU92bJDBLGr9aBH6IhySvI5f2BqV15bnIUYyS6YXfKu+BNBVxJf17iFaTURbq2i+giBHnAx4
CMRlc3N2VL0uXwul6anLX0uzmpSPzUx2QUNK0GXoSzOhuEd5i1fhg4d9udhvnIRVzvAVYxSDP9YT
0mplt1Grq3Ek904JBzWPy57r0e+klWFRA+3M9UlyfvM1ox0AlWcW25sRE3kAPxkq2kfYEtwjM9ia
EYLx0tloETEP/Kn0l4UvER2HuAXvjhHBJCwQf8m1bS0/+uU2pi/GA+DkT9AKz1TmNTuII6CizD1v
qgR+RjZ9+ZgLGQrzS54urW7u664kNCzGo0aIhnqo/lGhbRP1StdBBmnSlmxiJacq9gOuSvP3nkd/
KEWWaSnKlx1rc//ZyzuzpUp40RLbTduchT4yK4tRh9T0FA7WghlaDX/06PKsyIQmSP5NX95c/RXl
DGPlY26HesiUtDq4Um6lgVddMjtz0i3MM32Y9+RTfTKQDTmzIERxhYHyK8z4YH7mEW6NaOoar9Tj
Ysgz3q9zhBbBPJU7REZp0AFb3C5LCeXqZ+t0MmGEtHQubyuXV1Ffl+qfzX9IKHtCsPSbo2Sy7f+5
NfH1iGAR/HSifpBhxH99BwBwZHKVHYONp0fr3yPIneeZYoXCKchqPU+gwSGUZC6gQ13CIabSi/10
/bZ+t71YbW4oFPF3no1XRcBowNn4yGDJICFJ5AC4RiInhv6Jz4zG6/bOVpOLgOV2jTKDsIf/c7X2
nwU1NMIW8z9maK+/KXXhv14fbnMyvj3UThdqXQXslXPUg0P8Yx5bgdzc+SpFKa+Q3qTyzoFVks7D
fVV4i7ZFRXX+/+BDEJ37d57SqEoDFIt1u4r5hmjNqDCJnRx1uz5yZe6hd31Tbjv1lJAR6te4OkfJ
gdKtOoh+d0OncWJzqyJXSwp/x0fYB6lpCt+J7F7eJ6g0ecsDCsIHT5SI7DkMNjU/2s7XDWO0ybE+
R7GjNcMnYfnxCc+heSuP6rtHReusSF/7BM/sMfbIXWVObSfpTE4lZF1R1X4zUI89gj3NH5Ev2qEL
3a9FgfeEvLQ6Z6k7Y9k4I8/8ccIwRg0jAQfgfdlEWYd2gq01vD1A/Nd7n+cP7IO7UeIXIuYfxEVe
o0kZUllko6qTaoy39xuF+SLy/2FCLGeukmE1u8GzTU76g1k7REvfM2ts8+O+kuFQbKKIaJvT+m9N
NRhS0bB6gZ6f2mX4KGqdPNg5+DAbzbn87PGV8Bcr1oKaIzsmi3BCX9hDf53Dkm3rxSl1ir+Msn5q
t0IOOYwz+wonSy3hJRVRaFCwkjPgRKkqrBhCs6sae7makv1Krn/66r6032mbTS+ajDNoyEMzYiI3
TsWZffKr91WMStwoLssN2gQPkJEtKaTigOo7ao8yA+nWHNyN7gGmZdYHNKI+Vlc9QMG/B1c9kVUv
Rg21t4idNDloEDa8+4gAlvXMCwF+ljoOhBfa4ArdfN3zNSD0dwXbnTAKlKC0j7ET/Zb7E+Qv1E7K
r1HdFYAVMUHKB1wyDApmSRjqabVsaTeHO85vapj4faPUMZy+xJE0W4TjtiqMbXDN41eD7EBBbWXJ
kPiE9FFkKoG5KAac1xjYgwCwTvgRKYlIigJSRp79NYHtKa2n34Zy039aQXS+TBMPUO2vaxm7VkT9
o88fUylA+myLP7YqNgPJbrrRT6hZW+3JsNRb9fpE4eCWWcVlg+It5s07bOLzosT/VtswIuS1jjO1
bv2wKOcrRyg3lDWrWIvy/pvIzlSuF/wIX7oBndb0ufWraOVKUkQFuTX7t/UZa9MFZ2izb10G/7Kf
JB1nH8xPDsDK6pVELru2rGB+sNi7MQpaJrF/m+DVUpZPnufS81vkrUBqnnFEuVkWpb1FvgGmxV6M
CabR8gOFFQXLmGsJjscZhRMvRjz3BBYc5idpdhxKZSsPSERyZ2sxHDbUoOG2In1VA2ivSXs3Zrq+
w0xwhWSn1PyxtNQAALDPOLK/nR7zaiKd9FAWEZy/SvbZuzU6ri8ZPh+LAOlAxgxSbln4bRS1ZQZZ
Vpd+I85r/QNOqgI5Qzs21tHOrAQ/srXMePZmEcXkqB9bs7lJoEipyg84dX/LRYD/E9frW5kO11Kj
8OVyxBAQMALk3JsDItijw7eqMQO/uKQwD+8tlTp8vpFSmT5BWkMIF35N2FbGUUYHFZQGIQ7SjQ6Z
NDrYJKjN2xMktRql/3a7MtPDqZ2QkEdaMgBxYOZRHYLl/ggZJdlPDMtzjHku6uBEw9EEZqNODWBi
fL9bHR7uA11yEFKi+ueArF5m5zEQOkcgIboabkpKFVsNvO/y1dLde3OkIkJZyiHI/vnhzFiYq6EZ
bTGcm1eIk9VF+cZyvQmiIzpmVXL9nsPTMz/vtuYVFRhEBuff9QLHOwLXM6Z5xaVoBffQZcFdIYGM
Nk75gu2RfZul+4bV9lVe10YzHIYqYriQKfOSSr2ysC3z1hqnYrpMFvjtRaaa/76RnJvtEDHk5vNU
ofUORI+qRIpDK7WG5Aqvip210tuO39ZGg0LX5TY1oHRkrc6rCuFQZwoCX9SfdC+z97kaCL6RK1VV
5S5Ojc2prX/HtrnLGvfPUyqY47uBNpYpU9KXLSF9ba87vl4WiY+ZXe+v0slTEjRZWRWw/SnIYCt8
DQ90lOpurZOsIkqIiaAn3pLBiuhPE79GSCpxkCD6DYnQE6u+5U7xrnEQ5DA3PsXrv4Ig7+C/7As7
0IAAMEiLIvNhcAS4QTqF8oB3qefVfnGL5GliLzs0OgNInRqbsK+OdjXMFMDhB13KnckuZmkir853
xoGa4kyypOEJY7NNpuj0GSKzIIe94cmywU9MQVZ4x08MBmhfK592XS2Y6umYRsYddf9erBQiuhD8
GJeWtjZy9HgsgtHc31sPxVuAdfdbSuh0STeV1JGQFd36QN3HLGI2nJeFOr344Rgzqi9lHHON0OjM
ruwCpOVG77g5qQrAyGdnzjw2WQiJxdtttcXRX7lGYZWjYyUHtwOIsVWxm/7gM6LHLWEw2jmrMuUZ
vtUmZ+zLCFgulLQmnxAXnX8nNETgIZVHAZCcyjaLm1okrskqHisROiouBzWejEwQg58KfULR847A
HqyECZKCxCHVVFriaJNeXQK1xGDjB0v8+H8k5bzKqTXbgEjY0i1KbxaZHN39nRjZiY+7mFZTDrMA
SMZMSnbMoMci/tCvkxOP6bPEJd8FEgfPa65WDKeUJvxcS5UBwiHc6VSq1IEYeJMj1Vg/g9fnv9KD
f4/uuSXqjB42135hxMRUc9rqDmfHU+j7mMtwp2yLognxI/3zbbYWXLiDbPDjm8ywoqFDFqwMdzD2
jarb4mcLIcF6UZJIqDG+9mf4cyU46jzW4aX5zf9BHF7PqFYKa/CR6u40EWHKMYG/K4e0XT0S+/Pr
Cs3ja4td8ylpIyOI7LPgkVNNiRTLzUsq43Iaynl2kzNJ5cvCGFg5ozc0x+/wxXp+uPHz3JixqnaN
63VIIPdNgUFMKnoQPLqRlYAy0YXn0NxepVFFms9fPb2ZmHC4Nl7jX7ESjWg10XvXO2cRnm0j+JhR
b3tTQJCfaamQKHFuwPXCysMX8AzLMNWHxB/dte2bS2D4eX1//AmSvOht/NS/cAMw82rlaYuKDeco
Ba91MSMmCHBLwqJXTXz7MUs5GeOu1k03azPkmQ4++O9hB3OnB+BlWqcCSNwMklmp1ZYpZSdLOdEY
qCdYIKEPEP4BZbvyD4Y7KY4sqvA1vwElc5A0oVfhtzxQZIg3GGoGNcbEQIbThRmvvKfQ4hdZLztV
eHQFD4LTka4Oujc83tGe/Td+saxwsoxQjGiu6xHXMpwYPbhkYl5pAJtTa5/c2xLU/NkoWYSFVk+5
DpIQP4Fek2sOROB0jyauoSvwNKQ7+o89TbaPf/hKJrrfO2+grQRVcWli6CgIwrzxdE8PJEIsKMOg
tycqU5zRx5HZBQretS43aoOh3CC8dToasF3qN7inr6wE6kvn77qYXpA02kLMJ51C8BCp34Jrzs2N
/o4V0gszbCRyy8RCnXTM6JuOJNy5uXfRv/PeoSpmCNesOa6aG8Omd2+/SjaHpUwTjkQKRciBufjC
dyCrSs2GvaN0FCzzH8X9IY9l4bi4DlxRRFAs1YcOmBUzX2UOgmmSpfsWmzzzVpBIJ8NC5aQwG6Vl
CepiGLTGp63twL+ZGTasxND7O7sG3yszB83kzT7ANUEDV8PELaBKH69A4Fpez6isupl+edfaVq5y
ZvUQe4uP9bXj3b5kqSXfWv1esU6wpLgn8C03W4W5b1d4HmhES3dIdJQcOnjJTvuSbYXlx61VYsJm
cG0UOISS0ruiGe2ayYtk2m/ah0DVEquVj9OF5mz52TlDrJRgyCfqr+gi8Qlnf7mvwsXMEmn8JXZD
ehL5UND0YU99Kf/PlJOHwd39NKczj0bTfpFTBBRW2hOHcr85qje2BACpwRzboseW/cbdoiBlZyPw
DV85/lhXa0HbDV2pQU0rw0OE03+xPaTdW049AcXFd0Q0yW0mNNjVT5DLOv76SXL0glo9pIUKXWT6
40G0+6BtCnLtD5MJnEee/fRcYOKHWGT0HP+7l19wjyoi6ea0cyPfPm6577l4QuRASnbnEjFO+KaG
baMr5CDrNcDdfPT7H2LPAkZTEfZKGYW0yu3I0xa/a4057VytPVxDUlir+q70PrPRyTXmBg3BQ7UE
i7qyvhC9n24UtMxHajHvXDBGkbV22oPh8ixDuTf30igIdP6igqW2ckdbvExwGKDnkdiKDpKapBdq
ExnDiFGU6HBIuDWBlfHXNnEAF7ItlsWNPJ7o8EZv3OTTUYrxGqKMI8CRMmk/CH66lsNBlaOa58Ht
qtIK3+nMjjrtbGIT5aMJXY072NZ0Af0HV5uEfFmIjxL9CH3kkOPoAgV7RtQRImsbKuOenr4zBd7E
UYMdV+q3feZtYEyy5Dl0yQWJqueX0I7LfUXXSRPJJBk49mMgqnA7KRG+1IpkIPMBc+UrTdkEGrbm
JKu7Gunx5/2+MuZqc9sbucunqNhHarlKH8+bwCPgLu9coySdpxdmqelOihfM0k1DgbLoBDP9c6Mx
fe+yMmnL7XeoeDLE8Ws9krTWJc7ZYmJV0/4xnMIoAqr94x47VClHz+nmH8NSdIqdUsrwwdHQ9sdB
2QC+OT87vi3SpbefkOUv5S/XT9DBjLL0yIRigL1rKDDnEfKOnuJqtAF8EPb+e7S1O0SfqufHAybM
On5UJuwPfXsrIfryhXcMhrnfb2cADKE8sqop/4l2/vdEoVXo134dHUa75lSV5tz6dxeUBU4rVCyT
cUs+C7gCeFGR4xJeCH5zWjbZszi+/O6WOa+93lvYb1ZIyhscVMS3PxfJj0TBBo3Q5ZIGMOzkR4s/
WLw2lcZDf/bciTJPgwt1AFnSaW/keZW6p/33b3U48of9Io4xO+tKVqtjqY/EhO/jGKuEximyMDyZ
kO8rscO8GV8weT9XEm1Ptet6eWRbmD4OiVzO3UDlY/ICtm18OhyJvBhmu3YhRpnQ1Qq+79rQyKie
mN2ae6rCCfpkof78/Ivl0gPpWj9MJqv5yq7ZTDF+NOe4Of1plURFanjenzd4GNLtFjAMZMxiKZoH
m41G6gEFKLos4AcAz2FncJmxTn6LuZ7hE0v0EAzO23qemFamCVvXaq2zJcHcZSBy6rlTljCev2l/
3aGgL8KYQZniuTE2U7oYb9ogRqbZvFO6tgIL2pXS3ko7hbolN/GWItHX4zohKh8sSoj/V06BxWb3
F6U14NS6prClJkXw5DM56DLws95NqwBCJzGuaAoUs+QpA0RBQYansIAdRSI45roaQ//JAz+hTUp9
iB940JCxC3DuRezfdKGAcfSMebbcY5gHyO7xU0xi4as81gK+1hmR05TTHClDhRokcbi3H5sx2B7K
hXpRINzUExwNc/n1AbWcEzJiDgrBk4grwXZ9WrbSgR73stIphW4olDMbyBZeXY0ITP+Q+z6sXu/9
6R1XhwhXYZvkz1JucYyoeI8X/P+ocrgc8lBfvxTnuc0F6ow/DqfwQ5ieoBEkYyMVV4AIcgs64g9b
OswJnK0N2apglr5DhjJt1/9Z6xv2YD9I01zUOlBW+YM6ca13MhVIRBxS/IZm2NCG/U7zwwiZ3VWO
t3u/T2uzKKUJWZxargO1vXxBhnBxLWcD+k7HqGITde2MLMXnqH0//21PtyDfSKNQzieu1I9x2DSw
u+5Ml/gbdqzoLD5l+Z8lOCUtDmsn7hljU9xYZM13wCYrtR3aSJkZDR2fdv6oU5KUmHFRnjO375bG
mp0+wHRXW0PW60OZOHRr6WBePsP9hC2rno7pZNJbXKg6ukHiM2cYPm45PlwCzu46t29xFY9O8WJU
NlcX5rrMrQBmfoxi9PLuFsRMyiP4Hd3ndz7hZtSgthvCjiKkFgzVcdmMR3lu5XktjHprY9VN4KxL
PcfL0KTMhvxh4A9VhZ3hz3SFSMZ+XAthJ+thh9HiOF3QqkdKFVa9zXomnXJhe8aII15jUXVQwJYc
Yslt9UihlPw6cKHFS7vBLNsg7Ze3YtouUviTnfwiHUBCJi+7XVWusFdpoTqtG3WUlQ4skD4A/1WT
GFtLMnLi8DrA3c0oHUUdIfsaUVAAghXVJ2goqd/dx+capoX7pmP96EXsBr+3xB+KaDeF4AuKa69x
S19XEaMuvkTFFxhwpSiO3/TUEegk8vcHV1em6ugQ67m4GESAaxObgfUWCDoNwUbL3Wdqs3EckjXR
rJ+mT5gIb4zfabMlAh1yevmRQ6beXWx3Ms+lJEPBgLRS3fBN+kdCtGwtGC9C5mtq0ZEtCOdGQn13
qzg0pL9XbC5ynOCzG3lFWrpnjiibZcUOKaUwgtC7k36HkqOABqU/nH0WKbf4/DyOwQZ3G0+IwgqF
2W+H6b1zoj9sWp2z7G/bOwDpFRq0+TqW5N8booDNrWCBCbVj89jnMHBtCZej2re6sJyvMdXp3Mw/
eGs1D2JxBtrMXYSJUmVCZsBtM/ezqWmebihmhmGs7qvZXecfwm1sKzVnNhH5Ayj6vTRgfknOf/yB
yGCnz3pddUj5S8XYlIH/JMGKfvBMh+dHQSdbttpPRn0cGlFaRFhPTbqqPMjipjdZjDKn2rXpErcG
ZQeXi8nDQddksu9v+tlPz+LcEiCl5km82XfF44m21vWyu1d4/ziWG7B824KWKQH8Qtl3aYaqcmex
Addn1b4gFqgV0kdtr40mlDMWBYHnGY0eLa+zMbzFRtpJiNi1sC6/2w4N+FMkE2lByxxvO6Jw1iYb
3W/TS8a1jb5ieFGwwWyj37k2lYc/MffyMbH2qTnd0eEgwTSkI0oYalircN8uco2A4GS5U6ArxlAi
awybK5pPEDIfnuJSNyLvLxUzTzZKpZ7WsPECctvqrzsBiCFPm+WzUuKhhD7+pp3JHiIu7YcY+CG8
U7ggwJBS12yRD0RtPgMtVBDYhWQg6zXL4/e8XMy8ObRRDiM6nbgYGgFjRyT9ND6vIVzLB7Y9THBf
HdG8/thUJq2g2E9dK+aDaFJsGKNKi+RQOA7cgIiXWU+5YxUGiSF0JyZpshVVeIlmPEXPSS4Cd+tz
5aYxlZX/FeA7j0zocMBsCoPc/1KmKRn/wZAwoiEV8ejDjCttDg/YTaQASTO4h6VNW94YafQE1J2n
YCVhgqQj85jvue2ODF/JDWwMsEW8tSd9Y/HOaRwViqVE+vSrhSJSiIxnYsMLpUCbLiWGotk7odFU
7mkUrMFwum3h51bDhISOhsqa5CFpcGMxqDqjAUdfRN8TcTMK5bbdqBe48V1gmgNuT64IllDWxXjn
mbKR4g2MfMg8zyZDNnHbb60ScV1Hz1XxprI5KOeJPAbxc/R5rs3LB5xUE2ET3d29MfDuHjXA0PL0
wa3uHFyRUuASnVqsta5NOQrBm6p9UywZi9r3aSbU907zoDykp1YzvFvnDnSn2lpGk60fASD8UGPt
xK1mrJtDTlfJ2HNUvobUtlQunO4u4BERgk7LLdqqdVstRhDBt4Ae6Y59/nCby4Xfw2ro2ZBpxTo2
A+4V2F8gAfykvJjzT+v772N694W/ezc6lPnyyuQ3FMB6UrdJoicOQSmSo5VW+/0l6kf5SdjbfjMd
7wS3KyNCxzvKmzW//3J/hm7QMOLLEBr4oiMJJTmU6lfAiWeImDWmJmf5YMCk/MukUGutDfP00q6e
z2PSkkm/G1/lSQQv5k2Y8Eh868TGliGJGln9UEsnjTY/+DRWA5InwdzTNj2SlBlvqO/O6yNmIyVQ
qVh5nNITvtNv5okeaAL44XH9IsLWJVfMM52YGOql+cMmL4Maql47qk5umP1PXwrZ/OL/ZZ0r3Q+n
zXkW5BAxbgbaz0XhB2plIH8+Zo8jNXanOUHldqVpmLOwX3TwTFkB+eC/wCNJLXn6To0pQMGl4etS
4nXpWPe8Nqm3XStnDAANoGOHbrQJ3jr9VFO+u5YLS9SxTMHuMjma1gVXPi4NieGiVpbi8Zjt7ZjS
q16wJ/ZGJz5S8M+D38qAsmi7epjfQETDUGxhSGBsKSsfhfTQd3KvcqfkVeeUcrpS9OU4PllCPDEk
7ZrAycFBjWS8HiwfGyB0RicH+yVvbNePTQJ+2TfWXQpxwpZwYU+qBxoK0ZM9Xgp1Gh1o99Z5POXt
WCKYX4r4g+FpIYE0h93zCPp7ACAvXv1VplvXqxrITgVsfTH0b73EYEoR4ApKmkqfsYFW50WFYpll
7+Qk4+hygXtsGR2YrahbwkueCtHlYy73nua31Lhoyx2V9lMsdyNjrLBw8HaEgdSKwjzTFPDrJGhj
kUQJZ3u/Ieag2Escoh/BEr4LmOZFIWf+xAx+TY2B0p+LVPvO7T2LYuSOypDX7BnlnXpbslWf1uZE
SqCOlXo1e+v5yX6WNgxZfKm+GjeRrHnt95W04pcrBfs8fRzdjMszjNGB+SqWTZr7YvjvQcEAbntR
mFstjlEoGh4DlXJZYqY3HcC9SdjnoylMuwkZ0MsYHH2oIfXGKtRkm1X1LYTTRfBF6NcQ++F3HbcL
+jiQEowxxxnLqnpb2bxbWP8cIbcRSm45TOYwdSQQ9b9il6u5/ForT7J/arfaGtmZoD/V4wBFte1L
7+m++OaZF7rI99aNsHkYv8DjgdoB307m/XashJn1jVdvMv1U+Im5xVHw67IWGVEc2c8NVucTdfhK
iCg8U7vcqmoilvLFhGGDGNMFK1xzudI1XTMBTG7wyEjJwp5zGlA7hmFEf14GRL4XNtgsYvxVMSu6
YzA3g8Eht30TJsgV7gmGK45Opm3oNdbB8ANeGnjTlesVNtc6K65Ygk54U/miRdWiUkSvpYvUvXbV
OfwTMesHISiRB9MoBZl3bmsxKI6DdgO4KF+bRkE1w7mVK3sld7GMmQQSQd32w4IPoMlluH3jhVPf
fY5z/MHuFqRAOsELVmUQsbMxuuNBuIPVoo1HS7uy/K9+f2umIwkPqA4yJeYhmmyHKGQXzDrXzdqm
1YVBybBqnbxjds03fv+p5XhEVsKOpZACIt1caL4ky9JZLkBwp2wSs1MirUqgP/BaaEAcQwT8dv2l
CY4gTyTFIaRzqCXEObN7MlpCTTk0HqcUl+b2S1jdn63DSxOTiPET0LOht4Q7WfhUGnvoH/lYgDY7
5HRJoNKZ7DV9fd4orDD/RDssSd4uAFXfCluPAsw/X7EkypiSA63S/Ksc5nN/esnylP0nzVYCTV5j
+GZCIYWOLpMJVGHmO1ULj37sRn6wT2Er5q0xd0iHuydgjjoS/0dtCVfkJHP7josoijtYeqobFnac
vMxWfMHNl4Oqh8uS+cSomCYn06F+xJeQnWX41m4UjsAZgcjUGXVTLM56+kK6/wmJiuzCSQlKDOxg
JYBTVQdMV9izugA+WIrUcIplofMGhINRbtuCA3imiBoTZGolu1FX6nEYJgYg4VDy4XnqXKotcOZ/
Va+XbuOA7ea7jntjinlfoXL0OBwN/M4aJ/JqZtt0OgP5GfCtFM/zANjCewesTBQH9NHxulrbqGfb
Ux6YamMXEJPSgtcxh6sWR3j31u1cfAqpQKZxUqAE5r3HLHzgsJIoIVkzl6LWdkJsQ3z5RWRnbrTC
AUFSBkUfqzX5Tl4/n0V+/Uo6GXqH1qUg03bd6AOtkNfKEClLNLALsUB+eG6YzQGFvmnUkIi4SBXo
cAFjtVgt5BVmXHmGtkDAXVLD5giJ9lnYQpzxdesC/55294hgv4bKHzQgNoBNBKvYv5TFuCKfixSX
XUFz5LirjNBWXcuoJecD3MZtFP3ihFNsggjHdk4TsH1sC4Kd8Wv3v+8cvrDezInSki9lLqOMWdWM
HeICJ/rG1NrNjdMddaEdSQ5/xFYbqSag+emhEnSnb9iHrmM9CXiDifEM8YTgc1KsYc3Vc/HHu0BF
EFkaIbjmk9FVcgkdxy6xF/0UYCfaf1tVDF9XoyynUrrjfsMbns3tLFSLJM7XpPxczRMOW0dI0lxT
GwW/qIpkCa0SDj1rGWTjTc4iVriKDwRR1/MzPsJK2G6xd0QNKg9LTXy2k0LUmPMXAt6BDyw4QSjr
up+/u4H97SEqzpUJQjIfShsnKCnRaVvReMLEBYi1IkpA/Gh9nG51rLdeqO8Bdza1i3pHyXwMd9tT
ERp6BsyPSWnD5C8f+uDgy6MQuzrhQOYBjIM7xh1nlGhqo5uGbtasZO3LHWrVb5Y2duhYrh/pHK1I
+2dF+pfuMTdrCWUH0RQ5qsmX7q+T5Z3Y4CiVeopQXZkwSEv60YCxPZvkL0lunG1VLXSsWomqA3we
6OqlzZFMyPU/HIjkcKlTKLojeXyBljZPw6S7IIvoJwYsTA11w7NdMmCoG+Qa+VGasx81xEeIHR4q
lHAecM2oy8ZII9kJHw4TG7I+OM1gjf7z+MEFcyn33PoTXcQiXtXwWnBCwhrTD/74iNlUsJjPp158
s0DoFgxcjCDbkqebY5q2NMSMQgwVXu/6Ovzm5HK53JsE07swv6gD8ig+vWmci9JCL+r4qJjcsIXW
MHm0VwSTh/eaaIXjM2JEmS914H8a7Qv3D13NaaEWXsZDCrXSZCW9egSX7PyrvSdZMICLqV1YOosq
saucIIJcyQs7l/KykhOm1oHkiN+vDBbZxygXImlDqIigiXR2p75K6ssZhHtL8JW17xLpgZs1jP6F
FzdjtFMuGBf7fUHpclkVZhiTRyQldHcz+zh5G90WU89ksBFRUIcEV+Mu3XnmX0H5IbL9dIoaGDSa
MMLj/X0kgVcxoHVc+tnwbvfTQ3AYXjNHALGJ40SQtlL2bRYNS0VVx6s4AfWJVTdehe6xoyzzcrsr
QJRM+DzsmFGpHy0BRZZBO1iqpTbn0utsaMUWplL9GYW6nFTI9Bw3J9mUbGS5VTNa5r6zvHIWIwnc
CAZhEhPNq8QzGeByQspOBghOVfoyKH9gMsCo5tDYnEcLI4b304iAsuHWZuXT2JCgKd5qc290T5gl
d61U8Wm8Yz/W9RelmcmVjPRe5meLRoxcUuPtV8i94HZoitCJBb0aDwXazQ+dM5qUmn2JVmVmFBgV
RaqwOZg87CLDTGyGu9kEQ14qk6KFAqEfpfaINHRJunyvE3CALy9BI9Ku06KpLtawqzPt1N+Z7B50
mGrKMbH5XH6a9wdpCgRHoDp2/HhC7yJPqHrNrTtgXaN/1ddiNduJWnMCgCaN6DbkrRot0Eq238wi
PdKKVbZhQqv2ORARpKTFLlYJCv8un+huNVGLeAlmaVLjyniFpU4s6IVeLEGONrLNzqJNCfWlcX3n
YdUdykgjqHw1LCdqhA1ipbkiRmPy4ioTpaJNcSnVL0v8wZRNARE/QyfECbUwHief57Vtjhptk+Le
r5we7uA9cmiGT5GJcpBuwjBECqQ5EzV0n6oLr4IvXW5MclHt7F4pC3yxrXRxjv8N/fKiIHi1NCWT
uCx7BkTXVAA1xpScjrAdFpKks3Lw0c6CibSonLXr+OM+Tggl2w6jwhTHP9IVK33b7XzUuRjONyUy
WrBojZckk0awhli2BP3FgyL+K+ei3k2nZawn5h99zsdpvYTyEB4R+5KLVx/up7TkFwLOarDPIMtQ
644QJHJBhR/sZ7I3/Qd6FIVn0PTCm8z9w+7NcrghYI4GoGnP2y3s8zyitGH+jhUgeeylU/TtOD/r
Rnd+CZ2m2auELd+/yP/fau81WYRE59r4ODYpcDMp4vNgcURynSTyyMeL6t91xUT5jqXVLpx1RdK5
mDfPa8gJZCHyM3IYINkqkcDE8j9GozS2C/o5q1SqwHaISm2qu1rUUtxChu2VlbRAC8JYGyekExh2
5krqsQmosbHcGnhJpMOyasC7zKGYgnDARCzgU8iLcHcBLU08PDJOxue6/zB9Vdyty2RWfktH8jge
Gs4X3MJ0RNXZdVqUGSJzIxnkrCILB9TbaOzOpu9y0QZ7dOIUnBqUineoMRhohCGPigm7sodZqdb0
FWJDDkW0VKmk5AJdBa9SffsrZoievGKBR+BFssCkyFA8D/Pc5xqOqo4/n8niUovh/zCzg6FB86gT
iqrSM/BpbQ/SiT0S2NdhK+h1P4tF7g3dmuTfoWSini0Zj5j2rPKmBX7+TcPuQKThAIDR/q76HSKV
fqZAB6sCrW0NcBUUmYNi1U0398pqYRRaSljA+YiblfzUi6pNCLFqOX1J4sFiRJxZSjp3Igcy4SUk
UZgzn7BevTXEGIr11sUGBvSiZKXPdfXYTlwIt8ygdraCiIdtwRNTy2Uz6Uo1KZx5u+6YP9hD24vj
nc/vqJfWlVflxjdCyanGkG26LAdmvm0XMi5noZSzIUAOVyd0LhzH/yDsc9Y28Yg2t3uNwlfgqLCX
hEOq5hb+JVyRsuftJ+SO92RK/835wy3z7fMJKVutm0tkjp9T7LiAAKEd2CjMtMIuPuymUWrol4rq
15hOXRe24YBn6/PL8yakwqWb+qMs6L3m/+XrBl1jVuBDjF784DNjyAgb8eQI4E+YIKVbRMV0fMZ4
wiZaGcHJ6InZ3CLnN4urJBfNwRGaM22D9HfFleWTdbpFjs/94Oy6+YX5o+3gYWEXCoVlX9bguONo
gaAJW6uIk7GnNeReHHBxLF3PDQYR7e/D5aal3wcS13ctnBM+8kUaA+4nKWOeMLKS/xzXlW/8gcsO
XaCx1yB9xxUrv7BRApPh9Q+TNVTGBHASajOQ5A3HOWr47RIZbrL3Rvr/quZLbRp11fG0PyGUauJi
8LukaVH3okJS9rE6+UASUZfQVJHmdeQsr7hiZQYfu93I8e//+uHel55Qr54E1yQFWTsNvHx2jqll
ob9nIeAxzOvfra7lVUWdoSEfdFyxk4m1cpMD5uZIdYX33IpoljNh0NifXCuzEEEtvgmVEIbW7//S
bYO4f+p4ZCMI846KkY5pxfgA0TrElKBe9B3J81mDm6x0biev3cM883ksGXUzbrcw99SiooWZkFeW
gyIaspA8WbOhskTyFr4Sze2hiADQ36Bf4N8A2s528v1SeWKgtXVmyN+YdIpalfHSapjB05XXmTve
ksW54ubN3phwW1NKbs1/b8Yw9SsZxK/c7CipcS29pGphzIT1cOnBoMQMvCu2Szz0oubsLWsIl24I
zatfOqdoPLHIlqrT2J3HdoPlZrTyVI3xLVWOvHLOr/k3Jnl8UAHGwYwCKs7uLmg57SX1BZzTcA31
K20pFXB7hHpRAXQWEzOIrSg7WlbSyfc6xiIoJ3A/8uw/SGTDEXPgD8mqefF+CdK94GVfhI+WB7Zv
IxycxOesLcC3oRSBsFjaSwRW00W4PhCfsdiHbk50UZ1avdosI3/E+JfPAevkqLPlQ7CXnOp8euoa
dlEZO3xfJdiFy9ZPRpQi7mjWEiGVTxHJYNZII3QLtbqMnPmRA2pS9HGwHzi807+syMKCl9GTrDfR
bmAW+tkGrZqWPES3HVyCmQyYs9CLLga8fK2KgNMby3ii76EUQy+4UcZAN1/VAnqNJqBOGFAo15i9
uX5qopNo6SnBsp/rzAxPA9i6QJ5xmBELl2s357QJ27gI8EEP2ZZjC4IhfCC9coo3HOwifvI6+BNI
xGqRyLvnVcts1a3EpcXbgABf5gGYiE899eYSl0URuEiOnylAMrmpvK6/gjuczvukm6ViK/0SV3eG
B4UE8PB4Y4wDF8wqZZZdGf/NFlTEEfkuKlRGA66Ij5+70w07GwoAl+websE6N4fDweaXOzJotUau
LKLwlciu9gu0uNFz6Yy6m28teSuLEPZBWwg2ZUTC0sHH+ADLV8GwFvFxGEmoFHdkM/CrU8YTPstK
wND1YnGjLMNT3ZU1ITDTdQhzTnHN6ORQ6LTKLqLk2LvhhLcTRmA0ijjRhFaScKaGsux9YLfuMDtb
OzU1Ps/48gHlnNXcYQTdKTzHEmWEwecLEnfnDs+PvE0WCcg5K/HpvsNxzUZZqBZghKPgJA+a4Gk4
B/Hey9YuzjrdLq4uTXUEROkUTl89fnzNhJfMdzcHwzc/a9XbRsKM1+vSW45FvTREjNM5D5Y19YRu
4bbGXn2nZshiN5OOh8K3qngMvRKhdyA5MowPxwIWjFFRSwpVI/Vs1eOLEKTcRRuqL62C2WAmICKp
orvgmO3Uv/khGKt58EQdXbAdE0YDxswCfqbbfb/x8DHfl8uw0jiRKQQzER/AIGdH4ZJVJWFCd++l
At8P5oGIfM3cvryj6332/AcLeFhDAPwl7myKS5/XGbIb0FWP6+ZE7W6ZBija1l9QJFaUxDsjjQNL
h0/D/0J5kBEixDWe/+LIwaf8+OP+eJ89HnKcoag6velrOOO9mXryAlP/6S/azpwErIzwxpvjjigM
h7DGJX6sOe/ffFvee+PV46TwnfHd63FlIXsA6OYO9n0xe/uqXCgsCXGkpBW7Vkxp8VmXN43LLTJu
H5a7FY7TFcKjEYrOcNwcbEG9mtV3camcQR7w5ZCy0LNtHAXCJiDKzWrD7vSlZNXb/8NXNBL4mFD6
sNU/NyuefaSxpmJmf7xLBpOxlwpN2yw9I2iFXBgWgm4Sn2n9Pcgc8Zw6K3JfVSpUehBQItn4ydvm
eZ4vY8rl7ziLCYZCU0vICooh8bF1tzg3DCEU1u01rsDbITzRZE3gYcZhXGTuGrYO9sgtOtkgKbIY
C567WVxy/F+NjRsD/UX8Sq2CHrYmqYtc0DonlQTv9VCq8g9v4ui8sqSjDp20Zs0k7rGgHe5ZVIv0
pSzXCdZfL+GKlSULC4CK2PDomJNZ5Du+IjPep3nIdJPxaqA8f5NmLxIzDfCQUZH4xFFymkGXPNjw
9w7WIEkp60t7NrnN7wdseqtAdTwZg3dSIVpiD4tGqXfCX/ywVizJie7avrSuP/us0iIurZxB38Q7
bIOlakiWfjTR0Hx8HYLqlw0qg5RyAQr6ztKwRV/f3DbzaHXuvmk7mWtwsN7vTjI9aYZVgIAJztA+
1bhmhEsaNg8Ky95NodRboSNkTGBxC+gIHS2Qg/9kbqxD5h2Fm8AXi9o9IdZ7hZY4ft65gsI/2nQL
7w1pRYNWKXnJ39ZlY4wvmgGRAlnhaKW1uFYLJFpf86s1FW+iyoyr5IM/3kpxSp+nUHGJ9GVOroZr
kocqwI72PvTU9nm8v4wIpwHKPUNRHqv2NtlggOMw6TKWB3kWd0965u/sGG+DYTRMjphyf9T8Hrax
qX/RpTM/7uwJiihjh5mEFBsXi+pirIOrTtYVmN+B/QFqpb9ugRil4u0Q+w7OjBRfqUpT8RPpbJCR
Bs8VV7RmqY4Ja0h6gRX+fYvToInPBT/HfGChPQhiEnEKnZvUlCLEnJ3s7bvk+B17gEw92Zgc5CEn
chINQlbDwWoDfmSxdDMe8+Ipms4g4xPk3evhs+LGHLFkkQLUilJaL9wxljxHHJKLo6xEinYjk3kR
RUYYsM+PdBECQkL2LRw7+fLf2xOcJQrddQezEWtvwtfbfDBnbZdUghHQLGInB8wKGszo4OFnnRRk
S4ROOFRvnHtxSHcQtArPfFPWOlEHqhoU6zGFGuiPEUBNW4opeWuPLzvJLXZwS2O1zcDXiJxeKHxk
eFewixp/FrnCgfr4rgU1C0I4t5CO++6kS41Q3c/gQD7UJeFYNW0sqNUWRsB7g7NJucOJR0nmI3iC
FJMdW1H9xGABfVDfnGe1x3iqJ51SVBXYrdz9WLDweA8DGw0/+4RA303BxUVJRmsmdIcDD3FWR1WM
pICIbW95pPwfW6Vc6E9xKw/Kh8/MB+nH/GRUlyfyYm1oML7m1l+UrQnS0l2XhAQWSBRsBWJlvlZX
/Isj5RxFdVtgU1lJwscMM81ZN2MsbCWXGHH6f7wPmJkMlACGwXdYtWgYrO1qKee6w2pUs4a91qaL
6qBKObwA0EWQgV98RGqjERYIDbuHdB/PLfQYFRUTAD5IoNT94k222fYyxSQNuBRYGVeHFv8BLnQt
DvjSW6CGxzpxTQYCMt3zsoQMtobZ8JKPCrcMtubeFn0HL0JvLK8WP5CvhyUn8rnDFobdCGGKTtiD
jZrGLfSHUHMe0DIQ+AzxVDVWbe7H4FJANRkTzalcs0o7mdtoYsERoq8uRfVhHfmpYnRkdVOjo70f
PjssnoYonFk6pgT/PCjY3UGpT8njgPMqK093vr8sLSHZBJaZM/Tk2iIaGBw3fLC083a9L+L+/UCx
equ5ohKddupNbF93yA1MbtGp2jkV6VU6zwkK9saKTxdWicQ+UoujdBXiaH2Nc+U46UaWveDYczof
Qa5ggaP5wljfLLzNbgxnRK+bMg4Xqpq28YvJivgvWlr6E1xI4ARZgFf5X+fhFeAywTpumSRmc0h+
Tcd4Po1aea3qL+j7NfHkr52dwsG8dLMQiAQbpNpgU7Qbux0EfgDC2eBMdKrxi7FaDaQWfLiEjFAn
VJLY+jA76nLuMNpYYrvi5K8p7Ioh6c/j8oUT6hr3FNh+VP3V+pOUIJtjK7/eCw0eNoylEqoCf7BL
RG7GO1heqOfVF6S4Zsmva4w9Lb/T5DOjmkkfenLN0p/2pLgnj6O2BJrWUcoSF6mARwwuVR3j81Tv
QG4KKzRZSd5vZlMpU26+juKprYnqc+s/KLn1uwETFDW3+JfO5DZRADC0LmWZrr7JTEZULG/rBS/U
fDo7zHNURBzBP/1Ld5AzzD7Zv6OcavRnCOaDuBWQym5glmEFYJcmjOtYq/NhERaTFHxz3BNfTF4U
MnFGQQFIocsHD8NLbtMSXmHwLIzMFLO7LNDSaPe2ezJ3AYu/Ylus4p939kmHMVR6IGOS3xG0Y+d/
zdt93iLenf2PKeyCgPMWa2nGiHAGJVpDGiC7mGDfLtv/2MnLuEY3gANuuYVCbl404EydqvhbqZG5
ldcNziUOn7e/CUg2f0PcOumfSjRfu2xn6oMaftEk2FXQXzysZAkz3/A0BLKV+VTxhnchgqrPJbcw
wZteHGBrNdjcnf3015+ssN68ZDfIEnXfkiIuidWWEXFcRCM4VPOiYew1+IONknLw1SoagVV31lWG
BRv3WXhZZdYcFGx2Q27o+CFf/BqEpp/PufdTBCb2HbjtkF1UiBSdM7VLdp5QOlNZO4Gg0QXviO0J
CqX4lRU4Od43xzCKKlvpua4CeEEx98N3gmVFFz1ieHxaY/9enT8SRF6/6hKiqCWSQnlrf4WdY8bl
ySlBfklQ9d9aAfY3pPZ730opzaeeItW5rZ98BsMA86Fn6FPqe8cbqEfxkmo9G6k3+gDLhEsS8DIE
43zeropNfwXDb349Bc2ieaU6asi1OguRs8YN4H5P/wtwY8o7kAz+fDeWsAmU8pWP7bnZVe9GDgMc
ZelRkpS4rhQYVIpSKExOfaU5PZU28/si1prvxaBfxwbsx+a6VbI7Ge6JJY8yQI83sxfYwQf2GQHM
MEnPecPSEEOCSFuG3J3U/A+uWcL9zKwA80XITB/FcOpedBrcH4TQIC1FgFJx89GA/Ak5A6ZKxP0S
cxARcSSDXuxkezhPl0f3GUcDsKtjNqyIT/e9JntqIyyICwcfpsMiYJpYgw/Tk2J853PdiG3gcqYU
KoL55z6f2HouhUjUSIt37Q3Fd7MDzvuOIa7Qp0UWeQR1LFZ1rT6ffe5AZnL1rJ7/NEr5G8ei59er
qBXoOwvYWtQcjGa0LftzC4od33XOxVYKNEmBYC3wfjSkWoE4HONhMzBQHI020LuKxFe0VGJRExYl
hOrtcyKl9g4BVHzIE8AVoJWK1KJPr0YFb3nl5I7irJLJba/1tlBPeaHtBNfGk9qpnyz35fyUGzqW
qIIGtyG+cWMh7UJh0pD5aL+/UkbaRFkBFcHPo/dXxTumrBlxBq8cx28FBewwvTNEZE+xAVtfxPsV
QW1HoFbwaXXXq6bTN0y3Kga5mGaDcq6paerjnm713i05dCLidI+x0bby3OQPob4MvT8SO5eFEJnA
imetJ0OKQqJ6hpS0TvLAEzdyrDCOC+eIGHTkf82uDYdO7/yjjvCXZLjSq2D+eqUpZaa3hTfYj95w
Ibg3RsFqLS1Cf0t8h+WfkAVuiR0UVmpba/przZ/Ip0P78igN8wD1/UE2ZYcqnqUKZRbocaeifDaD
L7IDDTCYPXpRuF871UjfIzrRM2SROQ2KrBt4OjDbUoISaatFGN97XduGmmx4S9Nz0HCAYXN8ufSM
2J3G1SGHOI74WeZlbxhMbAzImfBm1DfNxKaXOP2GpAWRWKa9eHDZuetvHkfnVKysHfGED5NF5WAV
XSuJdAAWStiq/SKZjG+jRL4/8LYqiUpRCW5vSQCctBF4RJn0BfNmHMeqUKyrFmLoG8404AyuuEPD
kdA2kAiGYvDayXzI9kewmDsEIPUmiC9K7NngTPGesIGPv3QTZhR0y+FSYxFXDDps1wtydQpjX1YY
nwvohEWmHOB5hTiQukIDMib/6pKoTBgeo5Nu1wKMYO5pheL8sTAH1zRmgF18HYastLatvtEszPpY
7l8JmF6DRbB4HFcU6BYIhMdiqIvTtx7aj5sETjUGrsgDczk/84hSgUCXqMr5tFxMngFxRPJ2jskf
l4UwZASibwN8WMAzlgKwPBzYzhO9DfX0xXjHtPriyDHsaT5cClA4x579DO9L/AM+XOaNUPntcPIg
oYQJjKav40I841tBvSGIzpW0XxJRzFUCHLQNKvXNpo70/DPkVAkGZf9TzXoFgcbdfpF8Vat396ow
feFRAnUZKMRkA6EyoqgLQyLSoMTKEj/ZRYgq8STKkxBJ4wHg2d/7YaiRVO58mMlYVBmQq8j5Lthy
tNkhjQi1C5BgUB9EU6TwWvZIZFgDhr/Yj6m1rL99Oi60J0qYB4+oQTgRxcpGfBpCf3LwzBiyj/I0
Gq/wNPo+cZ2xdCuJhpyoqfWtZ3LoTeL6yG9HfDpF7QuqYT/NbHb60jHigPdnehGIeVmg7XDAdVxr
GZydVmOo7Z5LgJ2W5xkCq8bwajRwnN+kUSpAWygpdRDgnVSgiSVnilwe+EjBTGklHkFD5zCKN+Md
bEjc9nzxkOLVRdx5MNReVKLyyUpOJc193t1iG1smQgz9DrOYCTdincu6ve9RiiVwroL6jA36808q
SPL1662LQHaCCrX/1FolWtWnfqI5hq1NJZydH0gDq6zY/7ML2a2FyJPWOPPvZc3Jbz/taqIHv41G
lTQN1XJS4KG9YoxdPYsF0Oda6Sc9vQeDMj+PKqiFgA5S+ytdnZT3JVu5HMCMKPmY8aWYM80HWUqL
mVQDnosA6k1ymv3IqN0mls9PrHlys2uNQRRlDTdJSEyLeZa+yi54Kyd4mNxQkYLj/ICSdTeHPI3c
o7ab+BdTqaM7LCUjxioagGIWNEJTmT395qxCeHTO7feAqzIwlWMl6IPMaBOAnd8GrkAsch+U0hUx
fLBgPmsWxoUw7fS5z9rT1afJIb+wtjij6UeJloy+McK3rLXFnDv4mBLYsF5vFeO/ZGTZqig213Rs
HzAjfKKZYRQ9UajZQxDgLtNVrkNHNDduDqnze2Aud97/bb3NeMskVbLiQvjzzS81AAk3Kz6XoH8z
so8IvBz+f7m8gYAMGZDlcJwGoNHXPoE6H1p+Os3kC0eqGG2MtRNQKi34Lr+4ZVP80bzD+1d8bObH
x5281oOdQBbt82fiIA4Q1hWdyzA+V6AFDrHeqFKlFoszGsYUyJ1K6vlkqRiE2AThJN3jldOlogeE
Mgy2LnvRr42vt42ojuB6Q8STlS99lfkBlAn7JK5HPzpEdag4Hek3Rypiwys9upZXNf4EU9YRRTCb
3idWht1Heg1Kh9oWgkk3xqmSJ9updk6TZSXFryAh5V+Eu4Uon9CZdawTSsYBe1CvapwoE6da80YG
e8bhmJmzT3k+/Hdb3qycMcpP5NoDLjJUnNF33bjXB/ZbY1VctAQAYKoIDqqYXBa9Rj7A8cgAbtsk
lf4JX8wDFt/R5nLgr7/v5x9R8QWr6lyvuR2Cqrn19siaCLBXb7GfF8GD6FQDOaQY3KNvSmyHJ7y5
08pV6HaiBQ0pBw44xuTzb0hYUeTjhHI65J0bnPxR0brnvHJOMpC0+V+k/05flAAcuRLpmq1mBCA/
7hdp/vlwFw1721WTdWoLhDdbt8N1KavrZfCMwRqagHXqtzXxZh+xIqOl23VXwxZI99gTbUCLq5hE
vraI7UK3Ari2I+cEZK2VcXLpRa6lsA1jrPOBLfD6oH4xVLHVpId71DVBPtgnkjLg4pnBKngBgxhN
eEAJCvW2uLpbhZFc78vHbrybNP1PbGHDuw3DAMgdafMxe9XZ2N+VKdiQgHd/VpB8LOJDGI7kGanV
pHRCZlT+yIJXn62Cu/lVCtpzdu5cZUZgfXXSdxF+6ndadb+3fh9lc9IJ46NbZA6bt+wva70Dis1S
NhrXT8wiZF97KG75ZkQtKq+WQ9NV2B96mDgGRdMRAZTa6ONfYA65XSmENuGqAX/Puoyb5z5ZKY4S
lX4doUxLhRe8wf1+OkHbX5ZKnGUcPAua2s1wc2REPuQ72SNsybBY2bJcGpNppc9njCRmOLjxJ5Dj
e64TgisyCGnLqEGcqH+eqpbY7MX1XA42Xpa5IiVHtR9npXdVIEBTHA1HkUJMo7LqFF6/XP/Mptmm
6FEitvaV47/f5x1/SG3wFAGoEyLiAoXHocnm85QPY2ZOC/gIM9PL9c6T+ZIP5vhALhg3OegzjBDd
P6IJi4+K0UEDh5ve8mr4wT5z+i7Z0CueYjOdBhzsN7LLhwnHR8wdEOrx527bWGSz1Gw2gz3SQPui
v4ctLPbSE9SstYAzkaqVH69I0NbzmK80xUeAQNlnJ2RPk+rogdqWPC/ULKQ4KaHxNnvOGfLSQjwE
bUU6HCtM6OWJsHzGG6lxbjWg5L/UMs5B15k9z64NTm0QOBVUlSvAWhafj9JVMzjaJR3oVB+Pl6Ts
D/OAoKO2aLSs9KQ5YyiZmjnesgnU0smK8rBsMYw7KhBtG2Kwag5shhz6FTfgicf999ct7Y/oRIvs
tfewHpFwYd9fr5jnLt1ZYn2wPRZxlCse5tB4FqwRMOKuOoWFBcZdxymqI3vCglDx64ISW1VC+eRF
3yaTYSK+5I8KvllUVe1HcJN0/Msncw1udD9Pg4UybOeVAgxWgt2YUaYL/O9BmMcAfwY7UADeqqg0
SWT/PIQkJds1leHrOh9oibpHz66NSVfDxKKMB1V3ipQhaZaDI0w64hqzHio0lguvlqMbZMig9PJK
7E+S+H/BMrAUBD3RTVDVQN7jrU9HjYKGjJKMIZkQ9QkqHe0s/3buOTODGyadVkIJ8x4L1J6AoQig
BHxqYaAz8mRfX6c9C8MZvNfvv5VwEoQvRD5zTiyogp9364Ecf374PNsIhGlg2/lqtD9e4wjdSZyo
3YVUAS3VITBaX6vVyPCNuesa4CdYzt0dDRL+i8qzIl08nz+OR+IpIXeu7Ax36fEpnCZAYiqdyWXG
yIrZsZv+SxMXnU4fRA3LK36maArG711sXbtPapMSsvz3kTYFnFZ8SwLEDugU5haDaJPLDnFrBHl7
NUFTVMCdRWv6yURpUcN09gkxhTv82WBFkRqYV5IFVpho+VdEb5ymju9iLHYnsgS2vEuwiXb7Oup2
2Q0b6tIIXL895Nw2VApxISCIkHe5yuoTsusYz8OXFiLmYREh6z1ikrpLy45MhLl84KOMHQmet2H6
cXB2EHaUK8koJpsUr7VTjKBW2wB6pGLy6d6ydK5H8jFLyw7ss9HKkoy9fGwkNFD6bO78oDW59MdT
SEmTHECgDwfzZTURvd9++wv9kvhEHHnUPX2/qqBL548vKBTyRwvTgtXGYxLozrWIxG9sPEEpHZ/g
L+8WXrMM6Tshc0bSqEgDbvl4/kMVfsT+ZKexHpiQ+6Tz/0xAT7ol9IaglaOrbhChOk0iPz+RUBQ+
0Ppc/e0UE5HCsSjQjp3hadbJ/5xhalaCTHp1FWPk/E3cyhyOWQN1V2/Q8qi/5gWnOjzVlhuQ7cHF
8GQ/EGNdLG0UKAtSGSWx3NRBOjMvfwQ++lG43utDWnbYSvJdGYIUv0Er3AI9HeyF1zfpUCwmlCts
qxlYK+eCPZeANfOD0b8ZzeKJWtne1M+82opEXaL7OIDMsMUCe3RBfzZL3ttJHdwS6gwfowyqD5IA
EesKxSZKD+qADNVgDL8jD87HIOmaMhASxBwHh4XezK9NL+snY0JDsMUey8uKQkBteBwrMQUUsIAv
ZI36Wn5mpUY7XTEElzEtPS2q4+gsfjk6yXhvbiK4cVpdyi5dZ2EOJYNO2f0+QKNCSiU/81Co8kPK
SBO9fGHa5GCdkZX60CgAarWx7xFshUuBAEYpqvfWWAVV9h2AgQSPF6+HGwK+q8Fw8ByV8UXAOwVX
QI6jogqXuC8AP5h1FfDIuY9yUIYUrIPIOtCr8FIQJEkIS6WyFGAwk+ICQB7Fvc1QFt3UEYnB0Onu
E7d5oNVWWu0OGiElN3GEGFsEu2alJawN3SeBXSsME/JAZ9kBu1jROZGDllrWFcnZDKAQQ/1fV6vU
vMGEIQ7Td4HhCrz+auVWARhlmaUTP+uHg4nBflHVTZiA4sNFAKpzjY2BT7Ife5k52XuTmyZr7tHU
fZfknzXDM1i0jHNtyS8/uyctXSNvqFap+DNdkFM8pBzaYbFvnYsVlQbLmLW1aPRYlwmDDPpxtdLf
66UmABmnMU9cROokZ9RSV8H57sp/2vJU44kspn5E2qDoJD30R1Tf8JgBQai+YDc4ydluzyy7Vgov
hgnUpRNBk581PRQApfWh38n2akK9OFm6vgNXu3UM54l35hmts+Z9vWDLwOshoQ6FaBkQHnaXXUth
NJOzSvLZi2ynMEjBxkQPC/jfZgrF9THUlvTiQeMJHKf8uWlzzleSQTijXhngWgiYQ+auZ2Vtj5HI
0Fb0D3ATEhsZWy5/hBRzfYkAZX/T9kUnB4+v4Nr24u8sEFZLoT2fBv69zOpgRvpxWnQbS/DxyrOq
mabu7Tiwgp64YwjSLgzlXdPJsvtZoeEGNj2xeq7beUvsosCgVzS4ei42UemKUEdnesbktJRLDiD1
SfRPPou4xJW5gErrN4HsgKA+yZhX4l2rQXw2dk+1xmPPyRzYseu+Hwd7NoYcM6Kz2WYxabCHuEiP
Ad9/4T6k6OX33E4OHesxwUZAlwEXZt+cDBYy0mGO4U/KoRJeGwZiVf+kgZhn3Tx+yfYM0HPEKfsj
xqoLofMN/izIAb6/7PIdSX5F6+ep8oudM1atfArffKIWkOFiiy2fehDp7vPhlB0KkzMhDftNVDeS
WlWRfqtexM0G/SSZzHOAz7KPNskTpn2XO5jk8ZzW5zuhe0KepnEEXyudJs1D5O0qtOZgPUm2bsYF
I+GS8EHt49tZ10E9ZUjO2a4atoG5pN1rxtB+zS9uS2KiB7BO0SpuzmVIIFHHRRjax3MtREQO4ooz
ua6pB/niSMAtmwGib5i5fKk9D6r7vY+YkmuXc1ccFPppZ7l+p5xPzEgD5EhX/PzEDYTZNCbPT09Q
jP4IWx9ZGjifz2BDlnCtxloplRA27MD2NWGU8brWHURGonQCNHMWdLuBOvJVaAclFnppYqXWvcD8
KH0fvVDxBXKl547+70iEb6pX9sBCVWrX+s+rXnW4h60bczzzfVB9MLXdrCWE1ZirXcCAoS/2Uale
4e98FucYynw3KsSs6rT8kakjKS+hvXncYfK/6129LdVQAOyyqZeQpaxL6rYMGJFYFq00Tuu9B3n+
K/Gkr3jJrScp/Mz/SV1FxCjAH2TXSGeO8KJM7xf0LVtmgSXiq9kejnphDTpxajk0c7/FcmB55d5f
vFZxRAs2yqvYtevr00swq+Sc5fKO1xc3UyOqgZ+pvSfqzkF4g86cRQ0EWU2QDxTkQMs60gG2Pwvs
/c34fnREYXxr98BwJsUWzczD6qmDDUMcWVQNg1QvS8ioNP5g6EPTMEcr7siFSAeDETzi84VC7eaU
uezUfEjc17KJrmdZLtY4lUpilyYdyC8ExcHzNVjtGknGCU3mn2P3sBh4N6Cns1Nslbg3x2oTdWha
oGoKUTWbbn1IVkMlAhoDLzq/sJQUtr+tc4bh/D1Pc1G1YDMNvY1GDnLuehSel9C3KahwzTmQTl5o
hHzYl2fTKEQhidGKl4u6pb/bqzgkKs08DQ17wos68jZkgkF8CPugWFUEFynVaM2KaUnLIAX3RntG
o9LY5KSFSWEQ9aNRTBR08Yle7pFusHeVU5Qy36Ph+uvkpWLWhALxvra/JlE3hFl7nPEgD8L8G9Io
wXwyHLg2G13kb2ESNYspEAhjlhyYLU5c2xJou89S86XMCychCGrnzS1j0bRv/WFkGix+jpl4hePf
E2bp6OenDt+yYGbRQaHTVwInmTTkGC0JwCWlRQO2BBGbmz/jQ25+AL/eFNE8lpwrlUZyVcAmh5z4
j9tEPKb+tK1IwX8RJFbYEHUdsty+1q8GJev3jMqwc4Ovng7zhC5y/3CHk15oqAh2KvazFQns7Cbw
VaSvl5gKgN0GI3nZO+UtCHLa371u+9BG7hHI8J4pTe5R0kW/jWi1c5NTbqDDU/EpKF9/C+cVprEi
qvRQnKpzoIg44yHz8dTE8cbmVsPT4KRRlDiMalqpfN2HK0MY4E85B5+7/u2c7duFGNZaqfohAk8B
ybkPSs/fjGsv1PoLrUo4wCWwv83Knqz6SRoCSFcKfsbiqZOglfd7NpzBdiRXgPKH6eC4+Jqs7E70
ZozSZF6SlGmZm7vYDdY0X/LofNiW19gXluRMzKJKp2d3Rte4alS/AHv4sNBVblmnYLyyyzd4zIGR
hdo2oTJtkpxdQ5pwss6oFvmKBYmO3lWaSg3ohkRm/H1eksj1Ko4PYw8Eq6Wmupr/GxiUYtusLPum
AVgDvdekJouVgu2fySLoopIEMH3u2A/iuwpFbODGI1XrX+x6TfL9Lo8Lio5ho9b9Ztz1q5sf0wJh
o8yJCcxw/5rMR6s9XEoJ99IPNNcJhTeZnDbML65/Z6qtg/sXERjNwL/52oU6UUT60/PMyTu05/CK
MSK6ndXzs+ljhBbHfj6nCaxWsCFmUHXm43MTp+Sb3fD9pRv6uX0vjktY+3JVyHwd7MbrQtuLU/k1
m4r0xUWobqdh+K5ceKPsIUKfTVhIxxrkPBySXump2RYsZeD0bh5WlUoCGT4zp3MgJ3y6L8HfWEjR
VG4gmrgeB0dkNyWUx50uRNAmPxP+11Q/kua25OwL7cob5a7c39mTbwVtq6X26ZIPSKvdSAFSKnDm
JnpYxevjYXjZUpQDHd+dXkV3vYYYMaSVBbJivxbs8qbWBf05L0WgQBo0uZAfOFrsMTHzQvO6ajOa
Iu7KlwgLWcCzWu9b22v9NkQ7W96Jyn8408QofrJ4H+vj5x2/Z3kW4lLOfyUDnsBEMwNug6kriSJW
M+Iu/+Me+ND0rP0oCQw4Ng9MnvhSGTzmcQc0tQDn662Bb9zHU+FzBVgVjqK+C1xOLLupy5DBWaUA
Ys4WgOsLK1kntXxiIhm3OiyZaA/FRr29az2aYqjVwPefNLpmTYRhpH00zaJJutmOdE5n6yS8IAC9
ZWTGJ3U7CYjQnclTCGRm/ipmDuvCW9wOukMff9C8gB+V/1j/7y9gA+jSki2hMW1k0MmQKAh0QxNg
I/hV4H3458o7PozIhdOzp6Hp25V3HxUiOamIbDjAyPcMWdnTGbNZ6v9ZMHr5l5S5qvNKMvEx5CZr
f8+aZXtiKDXqkH05jtPy1wga9JesWfxL/6eg4GJ/12KJfI1TI2vFwF+WFdYbHUh9QW78BKmEq85q
Fgeil+po/092lzDNdGx+ZWlCeR8c15vUS2P7ghTGgB4KaPPxzurClkN/v8pN2TE/jV/L47J6OBED
ncoIpCZeWgVMzSq5yHszUt4jGlNuqlyiB4NaGHGe6kyqwWcV8fA99LC3wXEfK+qoIH3Fjwwu/7aw
Zw4QAtRzIEsWQsJuSa8zoGM3VHbvsL+PMInAaYqs2zjDwCRxHwXDhSD3la4koXCPT9eK8mBVTdna
+7tuzOJiERXeDHoHklyE/GxK+QNpm4NhMfFiWRkF4Rd+cNK1UuC3j2O0O6AqiOWMt637/aWvvYvf
E06Pxfa2Hw7Iri7MbjfSgjUFmL10EMO4aKkdILC3SLdTCr1tGtvlPh77tJHA/TYZnH8UYe2wFjbJ
5OlxmUVGqyF6JCFlcX1m3onrYksiCcajF1cGnJpOsbEGS9k63LmQTRteUt2UNx8ySDAO0cUhwSia
lI+bmyVGYE8Uf+ZXwOpDy+B8kzAk5RwaIjxJpNnzLsM3i/ZdMmMWUcGdHeF/w288AMEAfjzF40bZ
5mDmXxFG8fl8/bZq6yg6VSaFb+a8UyZX+DnMTd9TfGnpeJjatnz9hcUtXyo0bgJk4h0O6M3qHPD8
FQ3cAu5v34wwB9Od683UvVbC0LYIWv2/JuXOAeSwXMBFInvAY/0gIxo+DNHEx/YFFVZiaLSZKfIz
PEULJy+lH2OkDO9qxqYFdZEerxTVPiGMoGTjyiV8oXld58OoWN787jg44sAOG8BUv/R4d8EvXhE7
r/UsFf/FOfx3z9mFsqRI43RFI9l3g61AoX0H3LZEfrGOZWx6uvhMqIAc+DanQZEmCbDW8bHUTbU3
ZYZBKk/MSpuiJP8lzuA76bGguSn4YlELFRAh5lIQuLGmHVOoUzy0YyOWwxXsE+O39510gCz6Emhl
DpqZVRvh44izNUdjsAIgm2Y7z8SxKqhX/W/xM2e/98dKJZRnZ3mq1ysakpPOEHRdnGWZzzM89dCd
q/v7jH3SWNBPd46GK8nkYFbk/IzwwKPrF/7bPcFDducCmxFz+yuii8CfnMDci7oWKnT7jHrzkOWW
uviJ1xYKkESuZdBbh8jSMUJGS+oKZTIO5nCETfh8pZ0GHs4BPHjVU1qz664A3H39AhLowwcfrnpf
yr/t88Iio2PXMx7plvDzSJucSYEDmF34cQYZSPRgQnTRF7tQiQtyZQqX1K34NV2uFhQBgtxvWQwd
6DcG2GdmDuaTbsyEBSFrMUcsIdSx+wapPOLZcv024QNTqXvGjaqR6HkLYSeFt3tVCA2kPg9wq4Hd
k88AxCSi6HSIG70vWwUddk9b7WHYeC950jrAMLzG9/7nvreTtOvB4iRrmsFotk7O3kXR2Y2bSb8r
1/K8E3JfxSD4iuL3EFh3YNWWal1vQdD+AVGeUuQDFG49qGY6TxRVZwAJLbUCI1jrDEZlgrYeZuzB
gMAZb5Wj9BpEWwhK20Tf8rE9aARkBvlXDQK2LR4NetTU1SslkPDwDfxnlYeCHar/QsATG593bTa/
vPMqYLQrpE89yKfqZ9PpCAG9+190faySb4tlENIMmcL0rc+mF7xwl3PtyV8YkcVEMaCPWTzbBP9O
Cp2GbIFe3PptOblavvCWBOgK94o+/7PP67naEF3QPmZduz/30+9o/9sDsxTHOD738DrriY3eZ8Ag
rl6GicbOHwRhbjFGT2KPgzMl5nDdqMaUmIhdndJ2ZS7rqtkSBt/98p1e5WFbQFN/AifPex33CAzs
6dgsevi7/p/iWIctAK8fBFoAIO+jJJ9tQbcV02HA9DWcpzB7i3ClgpR7IU/GgNXSOYSKZy9sTKWT
ZGYW1vmJSLISfe6UibIVqsvgPyLjn2xhHKPFAGQNGAXLpUff37g0MMw8giivkT8l7r3lD+LD7ubU
6WhiGsbhJKlvCN7zz7pl1ndXx+GvScR0PEUnVRYPZTyJrgtvl1EtmcS9KZCPM0xihYDgh2NWj75X
Bxf1V+0oCfBUZUNESWCI0A0+jYLtTo+hkd3/gcsJB6w/1XPAQgDUTLqEE4mXSDMG8y/lxke+dK3L
IOy/IPhfBBMpWeMUDbGqB/+FxIkSeMxTUVv2Z9J+yi/J1WQX1x0K2ZTxmjnZaLWSN0lezEvmoAq1
iY0gZxRbz1NZU0PxoqQBulagsUg5AyG4J/Br3tUkvdBgVyCabaSBtwLUgITQAGm9awyuudUHT9Gf
9J3SVy8WMbVX5u7iNPahLP+8KWSuNrnOgq7hnJccphYMJS3Qd6wqLcvRMqh7oGidM5nUWNqxAy4f
NbknV4mCbxZkZCeIQE3pm7LwyRnsSKUEsHTinhJkk8yEhQShb7QLQadFnDPvayNfp4avlq3AYYdA
tDhl45np0Mroxk8M7OcjMX6N0DtaLBGrIwVo3yJo02KTc6OwDejjzEtUWaeGVwtWOu+R+JiKgAJb
ZQRL4wG0HrRRugw6z+BQ5KzVsgR5f3Ckw5NyTWlUKdMK2BNEJv+44DlVm1CZo9PlaYMl8EscTMaD
c6WartXXhbODFjs3ZnN130uxSy2t6pDnmErlDvIjHyD+P3tCm8R3l3xWj9xQtNpC9HdJU6stq0ZB
5arYPoVyKWGUgaqlxRTo+1rSVDi2p0USX5bKXKWp27lQLnx3HiLISl4RDUDjUbMTgs1pDj460xvb
E8W/FgF8z1smDcvFDP0B5VycECQ4Bq6OVJ/E/mrcDAeuzo1g0qKbu8zIqvtY/fQzXFSF8qww6J50
Owmqip3Ktz/JFxNr9xNvZEfP4hGMfrTM1pMqND91r4H4T8oJbsVVch5Kmr4jtebvGYlKR7pRdAhe
2Kr6iR0FVV4VT8+9DkPRtnqbMlVa4683caL//K+OB/dBw2tJJCwYnVwoQReu7c+yhquHYc6zRSdg
PatOW5rGInlVRm17itX/92Hg+Hntn0fnR1rjA+ZpdIn9sye7G3zg9vUu6cW7U9r1FmIlecybjQnG
nl3dl12/9PE/trtMaSzVIfg5Z4+GgsxUqttRD2bexpXss71C9hRwLZVpnSebXM0ml6BVxP68oHYL
MF5shernodYX9BGghvw58h71r16K0yn31ia66WtrQtP0NMBGzBtj5n6zoSR47o0Yer4szCyogBsH
ie/24hjpiaL3nDIEJSQlaEtVYLFwK8aj04LZYDHiJpZ/Zjr0MWsk+n9uFzwJ5bEP9BkFXUtRkRRl
C6keXfwMYUtTDEcOtweIrNnvwDu7EH/7cDQAgmZIKregtgqOzioEL7wQnlcoQuHl6OvpI+zLMy79
xhM/+Qj+Up9aRXn9mNAyKGNILFkCjCpRPWdV9PI0o9bpOmYwQHxTA76n+n7WcMGtrH36tJUoejXY
M5yxfcM44H+rP2DYiIoi/1ygNamHgoZfW3MrzL8w3cv1M50fJeUcEoX8MOD930ylDdsW3LcXYfz2
/5fxsWiWaQqTG/a2PzF+5VKHlrQQS3lzU1m5+utmewsoHbVX7g0ODcQI6WNxPfXbbik68ter3EJj
Mcac4T+hPYt6u+DXRyOJ5LmtpfsJbd6h9mmRp8SxXi34cCo7+2ZEv1jWKBKeiCcmsyTpPyL4ey38
ASzgFWTyDKllBr/aCZAOUp8gTD1UkBdhJzuLUX2wg2UBZ3TxKjJlSpB2CkAgtOBfXSoAZkQoFA9r
IpceJ5ByO5uz9yU+5TG9UI5KKP+Y/P1i74yYWp5nqw7POWtD8S7G36zHykDlg+lUE3tr5E6vs+Ws
U6Gx09I2anBhbd8Hq0VBZtotUkGlxjAjJ7v6VjYZa3vRAzfM+i9DH60qezNNyzHqiQTWAZmHG17R
RpbjPkQUQf/Jt8iRAB+37652Y/pVM4Jh1hdVTPVLjbJlFnJMFlFIEOwF/j1/+OkDX7gyT1evdbUj
aAjPm+LgVrG51J0/eihOGoScifgydGgnGTkHe8SyUn2dATwjK9DqQNzkrADvbQsSgHf/4FMHDVXd
CjOiiQCokvZk52PQ6NNZ3bnmzb20foZd+T2IozZ8L/NUkZcA2I/O1kHZmv3mel+9Mg/03pSoCE0C
1VS2dunj2yo/50szJZgM8JYEkyaZsCccveBBxaVIwvAeEct89DRTrJBYSM4y0lGbgbUNH9sHCLk+
iVOENgsSbhXWIEHYRHXcWhCzpJEhwG5/UPWiCSkg6+ZC1VB2kRqcdCZnkP0boHuQPSCfJANppYru
EAmJrl8h6jn9sh0CyJ+KaPJfpqaj1xyxjofCrXv16CCM4Bs4xdrqXmE6VaQ9wzIk6xpofSs3vWZd
PuxDvlqIq3jMia8PQ4CSD+euJzgOUbgn6gmS5MXySaTnUN2SSofMpAzmHr4Wk3kqnEpZlIlMoAdB
c8bC1j6Mq7YwmVWcp6n/ZntikRqSJzxpX+9uhd+diTl9Ddr/vRSj21xMeHQsn/LM3CmQXwnZDu6N
Cq1EF684E+qkGukA5Ua6kGh9ZS5skOlDi+Q2BPBL3pQb8ZJQekkRdbw02ACGko+J6mQyM838ItCm
zF2E98xcaA5iXs4/2US1Y6dJbkKPfxhKiZ95XcYjr7s/SFtBPRJ7gzQYiR2vgyfeKmneZ2w//rTJ
LOKPMpux9fi8vp3Fq2iWGWeKehZVYgfmZjN2a3iOleaZgWmi4AWwZIt9alimWtBsYREzbdHjuFrX
HIKxz0RhnIujfgmn1nESqL9EQMrk4GuH3ed9gTmA8GfQSUugNLeLnxV8QSoG6ys/DMO3hjJvxDbb
raijGPwJoAVC0ad7n8ZC2T7PyyQedgv6btcMZcz+pBg+uLszySiIg1G6eENDSy8aLocxUt6TVDq/
K3xR8vIxZtWReHPoW3fA9drm4+cnNXlbBkksGoi+dkXfXG8Utgi5T7LHZQ2LsMuUQTwbHYgCZ7eV
ED0vlE2LtFCVoFGZxRH0zQI/PQ07PgtY4YPfoj/kw0I8LsoNUS5bXXgLjT9ofZihvi2ExnLXcpiL
YLzs4AzPK1SrUGgnJWo3GrF1r3vnyhiQbk18v4RlKtEMOYAYI/3cy7gsK2I3fYvjm11MyOcC5AW1
vuxmbsmKRqP7L7twz5HyPM2sgGwiASTPyOxntSnK04GAFax+LPwlku9LkP/3bg9l939wf9ZGDILZ
0ry20TtWaYC5KYS0PWYlXn50BkUxMZuAPmYH/y2dUaILHTwd9NCZ6iQBefSncfwL5jZ/cm162E+L
OwsvykGCXEwpuaXjRHI9CSTXrB45hxvklG1W5dHx9n5F9gT9BBmQSZ3BQ0jHBMZ1Vwx16HRu2mBr
7IPCYdEIF3XpRAG3dTcYHX/qaaipt98IuXFDACJKk3i5ajeJKpC1/3vqxbsICHNdFrI6n5QZ1vq7
bcrRTspP4feOI0QfkGS7wcHDkxwaNJgXAWB/Tee9zOkVyLMQbPuB8+3vDgwsIabZ1W5O3F+jmajX
DWDnqjRD2NfxFfU5X2R7TMyyxSQU1jImjh7yVPeLazSK2ftKDIfC1IvlfwNi6RykdgDgTkbbYQPA
HvfHiif5ktYY0eieEAczx7G9R/1OR/CnKspyNuCp1R9qJmcA5rCKdUnNAoYxzbXwWuHuFiJaR3Sb
pWwQ7Ufa9GurPunDJWFPtP1sIelVn9Bdk03qllOn60zAD3lTH7xFsKYhlVHzI7mf0wPPp2QQuCXD
wlYDEUfJigMKioB5KxalwvIicnevxBO+A9KMqZ7bny3Y+CI6czpAkiCWtwcyjElYh7ZCYOupltVF
lGaZB/BSnJeTH/YpJYHH/gwe2qrzyJGlPt+VxE2HlzrBqy+90BgiTOLXg/D7BPKiNKrljWpd/PvL
545/TtQpdRw2NuEr+c8NrNT0tDAEfTNVKPG74cSzsA6tLNhjnE3bGIIi0ibCo9RhSwJLMAdd5R0s
Bt0kPu+hUm8FKrhwHLiIsRqrAIQzhJc8xg0neMKA/a3TzgVZ1EUm5R/MkC4Tya8XvF0GpvHrZ6gj
GKrT+Ri4ubY2Usl+t4gT16hz7jd0grYh2i2qSPWRgaO3dmZICZscSu3cZ6GyWDjEHb27QzL5R5ED
nChmpEcR8J3NGRXpfMssS7StzZFlzojVdprkYXonXEC48ZclH/VSAqQXoZ9a8OLZLwE4ymwmxgAU
W5qQBBr+yOp2jJrFHseJh2Hx/bpGEwFl3R4+zLTMQL873XBSdYoPHBTuvGjV8RkPqyRbdt/mgDgs
QqYNWencdm43npi/+kBgqovfd0ZQ07a0dnCfs3AngioyUYdoXL1R7LMv6NBWDezGx7yRu1e0ZrQV
+STdBWPCLkq0qskb2Pg11nM0hleJ2qXN0G8sD/lx837BtK/1WFo+r1W33kmV0JA0My07+UjkbQMH
rPb1YKQE3Bw6UG6YOszDJqQTKBybgftTjjJvpYtG/YEZM3jb+qbZchl8N4Y1PIQ4i/IIu+qWGaDa
CQjlbXASIw2VRBcGoCENWav2hJC24TMqxASzh08S6wiqjbrqTeE0N8270/x9A9mgIIexBpmQ/qLS
9LfHqWjjHvT6p2LRjHupA+s0ySw+yGqtPNzRG6VHFBTS+/mH60ZTp1MLQn7rh5q1ueyZbFI8bT+d
7bjV9E0eDaYJwE9hkhNlMIhQfcYMlQBiRbEhg4+hwsxzvbxiD4QpYxuQjdYrCW0GpX5h9IN4v7x3
2Bsq+YuGT5yvU2CORlc6kLN2yGuRyb9guvQbkZTusWjZqF337y5aKHJxHMxm6qJUtQKzCkA0EDSz
kM9IOj6vt3b2JcvTo6/nz/q3LT2c+9jM57hXJdLcAqb1mqb/2Wz8Xw5GOnPV1qMVcwyCtS+8T3il
miTZxdi3qnPOTlzenEYwVxiuILphN05tCp45bmPFgUd5AKgfBe6HNUt7XLPcDZ8JoAocH2Bb2lIZ
ZPm+1LEjfrjxJV2W17Q16oHGzA1LLitTxZtADXXEUwrV2BZak1iOYF08iH/g+r9eHiB39YVNAfw+
3PMfqm/zdXnIjKN/y7OnaRC1e9++9vrvKVRahBcQ8AVNEBtovCTLKItK/DuudYQcP3bCPKGmLwTV
mtbHeSUbhceiQ+1UvgutCtAEJqeQoGuKS6OeW+l6AKcZo9nrfh9XU8Tc0rZc8ijgumwMDFHLlbvw
0xcrawNVsB26+OP0BSNspZDqoaojEVhM5Rlic2U2BK406NgfWM7Unhz7r69Cu6DSGPb2zLozh0vD
9YW+rGPmrJ9r472DbbMnsL8GBEXP1mbTZm6b20QnI1XOXkpzzs/DsBFT5TE+cyll6bKY8/0JMAOj
D2y/plnqfWSoYvCAaUP7fCy1Nr9qOYCyrWa9nzUV1HjNoXbFGWjlusWm4i1r+xVERsXDkl/gSn4V
3WPbNvYwfoB2n6DdcyHzOz1HTOO19Oza1qYYF6AEPl70L7Y27L6tMbsNZLYey3ATj1BrJ2A85NXT
+/S0f4ywqPrqAOfB+bnDlocdbKtRE1kAuaqD5dcC1+6dcRl1bWn9npHs1fnDoPMxZxuQLuelykdy
i9CxEgaDv4cKSlt35pl2YREOz5Qa3ku4ryT9YWmO48lla/WO+YyxLuWGObAPM5TxG6b13V0kkAMC
BSPVKjQ+74V47JKWCLbeYnqEqcH6FiT0MF1HnnQj7ikAFX8vDCAax3656eQPJhDHLpfdFrxjV8dy
ITQIuso3uedw0bQibqdCmiBIJFzLCqOEoP+w0lqoEcopFUfYJKL1JH6/G/KxkDVui6okvUBuiVET
TwdK//nBsCcUh+NsVTvKGmQgvK3tBdKA3PVAVWegdtkRoQctYg/wc4dGTubYkWdxF5CkDfXyeisp
mKYM87x9qxP0ncY6C0jSb5Cd9DZt4SaPvCI9eWxZozElkYy2JEi1vgbQp/7WFEHXlCQ5e0FXNv+W
k3oTLSk0/rqPwoFsFwNktSMyrDyInj1LWpkvO5zoKnPqFFGsgN54l/Je/H/C+GDeiTDgKa6wi3uf
ritQ5xBybTYV16dOfPbcNb9hDR2ZPZO/vqxXf48jt1uxsnbPz6t9vL9+6Q66aOGwqZbbysl9xyQ7
YjP6SR6KLHQXhQRbYRtr753CkawVasP7CIKhqwEJ/RjUptWs03c6elNJRB/U4A4GAvtehOg+Lsif
BEjk6qLtgiagLMTqKFaG4RlFTYYzAm8Evje+iE/CMt60Vk0RrwQ5uW8Y5tYqRM+Qj05Yq6KPfCdm
tLvLpxSe0oN6fp3yavXUO5FCp9qdnXWN62xCG1BRAyOXfk0Wd8kEEFsuJCCxQnEcsJZEjBWrxkNE
uORbR/zbkVoyWnGcKW0NYGfmcplRVrQTZZknc7ZOhk8bBCFayJS1O14DGDXX6srEj1YzYGqGj5+j
GnbX6nUvQscVaFm2kCDaXcq+2Vk2JRw10wyrqibywiTgWcicZ60DetbM397OCmdIMelMQW7c3RFC
5v7/gRRgAzIZX+oHAHBuyZI7bquU0ZlPf93a7CnH8Lam1YfKVUu0Cv1clD4PA4UiovKX9aRxn2QY
LYG8fJe5RzVTVdgC2r65SZot5mx5SJb5QdkYVOg98kwFIsllyEq1wHEN21XopBVwJGVucVfOKx0U
o+wzHn9SZvWYx3NO7jRQqhwCQVp8nnTJmiMdCCCsy7+BjHniawKgh761DyI4fSB3HAwJ0lMG5xyu
M8esXn4MbF+aNybZslUyCs2NxAkPRJhSVCEt9HKV2r/RPmqL8KehRN341XVEJplePFX8b09bEf0i
MOaqyzOvmt47u0WO5VOIsjLROVT43qSUbwndYO9Mx4tME0JulROuYfJ4p3enX350Y5av1SZrNVx2
IvPMpwSpK8h2+B4UiPqOV/VPMgy68AI+ZZef39Wt9cuZd5595jDMz+/M6wqGO5NukvhhYzxaojZ7
Lk44cLbaAn3uGP0BobvjvvueqS6sPCu2IL7h7oUvG8ZS8B2XyfvQIbvOKmDETRcshso72mHuCgH6
/FUMX7SG6t8/AuUF9MaN4upPOVso16zr4fmhciO2ql9Xep40fhvRibUxqkVwz5K+q2BpXpWcMQc0
VXiTd7ck5cgseo0ErFZWPXjOzkT+dFh10WtdcNY1KbxK3oBkcy1N8ntcYo7uFSMKa5+utHd7J/yz
DvdnKIkidVGwkQ1XvRMSYeDFT8N1E5wLURzNmDhi66ScNJf5hMuIL0VfSnOAPFpAxmGmH6sq7cUn
IRF57RNrG2bMDTbinsNhuvsK7+3uW5v/0NUKkJDRnoEicv/IEyqhfJahMO/VcYWTDYAHVmvJcttJ
IjWK09ryFd4C8YokriF9pCr9PxBW3FBuFyEmyt+2NBa7rTZasQ4ZiTFGKUKHOu3ygjRydSaMQrmu
GCvenFVibKhfHfd2OXC6L5DeGyDVXDvbm8tdhiIgHjyQZGBC6L06oe38E0jQvAf/193sBJ0OuJBH
We2oyZzG9LTbRpWe9ED6mr/u7nZXF1T595IpQH/BGy691GLOyo/s8D1G73bkyaw0vKTVvw6ABwKm
fwqpo1+ycf6vb5gW4sSgUZmXASpAjGJJi8kIMVGgpEi+RunvUYatwI39CPdoxJd3Zxe1Y+rHZsk5
HJODHcsTlaIIlfWlJTqKn89k0kw73S8s4BEcoEiZlAg62WD0f4/vRDnkxYGW8F+2/OlSqx4XVD7L
GAjdB9DIjmwO90wHuTidgPXn4IyDMMMY698yJEpXzQ8nKFTqQiSpWQVidCb/LBG9xF8wQx5ARdGo
PXNQcg1+cjvq/r+/wfS0fSnqkm8v7GUBHX3HUruIp7mq08MlVuqh11npqFDXWXEAcv6ifPl65o7a
37WYDjwVR6Q5fdAtBa0KTQhHtLCwjyT04X3qzTBhvrq450wEpjTvvDrzf2O5N7QzPSnrgOyEIvaD
YgB8FPgSSGoU2sS96mbvwourYwvOHqCYchsyCrngqMsbLQ+kGVuGCo9/3DX4IHq2h1EsRbxZsVm7
8gV5Yrz+wOjSU8g0YxKL0t3YD6MEeiMNxfeM90tgWdz7LQMI/LMNbaXt6eN5tOncN4+g9uVFrtMn
VvWgJFwxlEQD4CzyHUgao6g6+WMVI5/0hvNcR6BHwZFrIy0dRo9uVHzRxC9sCJsXIXOzgPMUCL8a
d+gj+OpAyPq4Ly6lRpVDktepy8gcgwEOuhEzCZY0PULQMkPIYnfxT2sd1mmGKuumzd7sDrlaoLeW
T3bWHIbQmnKl7fiH4s3wsyfpvcfLaqA2ZYJQcHhKwutMRf8+ewEF/2LriLVs39PUtQIgoVHGBngD
29T66wXFAgq60Gr+K1yy4iew2e6h+SgNmKZ8ZiVJBycMpeuBy5DnqaQnnRfmEL6TN/nU0+ePI3TV
TMZrUn/0nUvVU+My7HyFrpw8ooE6anPQRDCtQdqiNBDzOubX3yphZHRSCuG3P4JMarD4+gNDeTML
J+lOSGQFoZg4nE0IpTuIF0hqPVyc7INdOJOHLlKmMr33u5btU/3AbZWyy2xKhEewoxEj60PgB7FC
Exl74tCk+TBrrX9hFW+Pl3UN7gxzVNxe9bwYiDMtRXSRnrlvgYUCd+81wJQ6KNfOyIaNrc4WSaQi
gYlZQWSe0OgMUjIXVz7pws5nZ9sHYzOBlySgUyTf0N/fwoqMaTre0GKe0eJ7TdiUfzYU0idGl4jq
1oFM+U2cuictvclzkFYJsjT+EF+AwFjDnSAm5RV2FPqjKSeKCfAbPYF8SDjY3a+nN5Pnlg5nicjk
LrDFtWp6+Lj4QRA5Aw+Wywn9lhZnpnnKsqE1FjQuOVmlqtU/AeP/Zhn3A+pM3M9pxRTe4ZpAO2Jz
Y46+NTN1HIqvE/foFFGcO+0CSnlJRgY43So4tGak6etR5NakuugvpOtSTiVDPsj9NEYtO/Kq4iFW
gAIKDdIrGX2f/FWcnn+gATFIiODD75Um14L46Y/zVTzHwG85DYWfoYQjZlNul35Hd6ArPexE+Dtw
x0Dcbqa5DHWDj4CHCrrazwhvMezmbXJYDu3sZ3FbQcV9nXsyw2UfXp7T5IW75ee4kCpPzH2Cj0Ew
xY3k/+t8zMpVszc0SYr03dATMZDw2MRcQjyZPOY91up+Gys17/M/bIFOCTZO6yNwOihLP2Ycup7I
LkzZFTyWr2NKmrzs+Vt1v31ZeK5Ouo3k+3F+ksEZCnd91MR1S8M+jYQy+tJfLcO9iM3bUOCnntIE
LXkJjBbAqKidjR1KurZZP9zRu5ekVOQYZR6jKmnnL4gVAv2zXn3SVkbElTjahSD+9RIVkvlhkOjt
fUFtVe+YtYbUuyH5jD9Iww11U0if0VOawUrefz8hPhrxE56EB+z5HKUW/5FINprqjx0nvLUVHVlX
0uxTKmHo05vLAZkGr0ukc7HrJcl82iJf+jmNBXc2o6w4nd5Ts4fUwasqyoAjZZs+RCj/sPnWuJL+
tCLkWW9HN0LCfZUZRF5L83Qqq7q8Zmm27Bi40V/DXCtLKuVvIwFx3zotszT3AHHmy4x8GDeU6/fT
icS8jPZ4zwi8M1e1UcnaaWETCLZrqCD+/USEZ56QBCT2uQdYzjfPEJeKx+iwCyZ8Le/8+vu9HEsX
4URSQCk+ohcsd16VB6sBxOj0W/WnZGVM0FviiuWSaXj138emRIX9NmaumRkhFISr+L0Yf+mb4GQh
2DzQCUMzVB7+1wFDffX0V/2PhIOnEcfPxsm/52sI89f/wlmNU44D4f1FxNs6Xt5nORfpu1xYvmHP
0Bi/ZqH7B2CGQGYgKEZTtq0f35SrXmKg1r49LNiehIVuQfKHHfl0UbAGWj846HIyw/LGIU9wIF91
C+6rQtl9/Lk4ariR8XFiKoonwV3GF+8lMO+CuXTmbQ3gu5oXEtsFZmxJublfF4ufi58UKCEbYsnD
+oVcz53GwYOv1UPYTofQvLLeRwq55B8Go65f1yvokJl1U9xtKhxEQOMCZ0kgNute7YY81BXAJ9Wk
oWfuwqs812DvWIWVZyRQFJNcHPlOwqA4WbkTm9r5etI3Lr7QptACczkUEyxFP1R02f609EDnpk2k
oo1H7RMsAQEv4nk16SvhpTTwGftK7r13bZQntZWcpiiXqFCaP/Z4nmGuJasyT8Wc7F4YcUZ45SME
cCI/IQRWvsi0FWeQorfHYJAPMblUkPZCs008PMV0Aq7sB1PAUMmT5ODa9wFlzqCW7He0UEwvvmyN
Rr3+kmAfHMw6fXegD5JMtxHI5WQXeRUAwM99mDbPBYkOzmLt1aFimtfyAILMe4P7KOIMLN4Uk84U
joxF0GpWBQFodLKyH8UHummSJzZ2DQ0QO/3v+u1JTFHwuMSwRgHwneQBvDQ8ZPxRPFihyrT6GlKa
dATP4UGXIC1SQLLXvlGpmSGof0Mofykq5b6SGhT34Ly0igHN0zTHIGSi/HafWMvdDi1x0SP7BBXq
04te5DfPYEUfij7S7unUIONAmFMwUArX4/aUAcI2lqPvQS+Snbaq4th8fFalOQaYspYu6gw+jNRc
hx5U1HMYjKxFv/Z3YpuuUM9ZAMPJtUzxLaWSTs6hoyUUj9v9dx4m5dzKDFHfu/ItQBSqc9OdkZIw
1tT6Fp96QobTKaeaH29r2KztNtZUq+WiN/nwli2HZ8q1jt7hfINVTX6u58goAd2ub7l0mbEa08pC
Qe1iONwEIH6fkHLoIGvId/A61msDCt2pu3tuMAfKzkib3CmivaF29OzvhdYOBHacSvUnKN74iFAd
d9DtdkQylOUOAARAWrunltL7ql9wbcDMlVhx6EvhqMv6cIKt8JFWyAo9IOs+tXk9qEkb6JV2h4Jg
wbDXmSXhrqoKQF4R7katHTa7Hdbt4uM3pwzNe1D+f6yJD5j0EbRKO5ySbz+u3g3tEss5CyR3w8qd
ihFyAJ6E8asXz+HOjcAT05bGdJOVdETEHDQvMv5QXr7650i/qfYC0n/KcEA7xjE5/h3gQZpSkuDe
GNmoDJH9KA6XxHIyTm0Iz2wMpIsxBfvxNJf9iOzX5X8qztlHTCiupkbR8/ncbN0fJcgcBVLD2vx2
10us++/DrGanaXdlf9RmnDtKTARA2ckjb4FJj+9JTeY+gJUdROSsVabjMp6jfQqU2b0+/DgyvZbN
i2sqTkPFlO0AOau6h4QbIQhg2yxvSnY+34zDhiLZ1YpvcxaSfsDKV5oNwrI3npIsdxg8w+rNROxK
zS3dZdRXq3tuZcBWDzRwazzOscccOj3VbT/iBbvygXo3LddgP4PG5XB6Puj2lIF6Oetu5R5a4MMe
pb5tV+7NAQ5x3UEUiPTEHj/gVJOGHF3fkKuhUaqxqrpKL/5UkL9iXUXuPZKh/hDze/Xnf0QZhl1n
xm7rPD15DL8o2plNp2NdUxo+SmLPRFuRIIqjZ7OyQe3jGvISEy9aHu+NKXvZmAF7bJrERw6R7Ozy
3JrMsv06IN1rsLXz/guOW00tZo/3lH/iACqwoLvpFBR5lgvxgcUItqympym+dOBMYX+bXNj81yZh
Whi+N8itByACg+qtdqo+rH/SCokhCWpw5NaZfJpXfby6SHSkC5PY2VmYy+E6kXxLTY6ePC2M9D6c
JEAIFfv55zmC52UYX8tFx86Uytyx3Jl8NSY/QQ3VxB3YtNvoZ+X7ECW6WWouUoGg1t4EQjBdAE1J
C7N2woWtG0CZpiFy8MQaYH8JonXOUYPdGuhaX9kqaqS4fyBZuJVef4ux2/xj0lkOYStsv1mA4nHG
8hBQwMNaxuCoTtbY3rQuumdbqAL5F0k7V4vhwQM599pgjo+JPlZFwR/A1pJ34HLBlyOd6M4xTmSl
iu2fosl5iVwdToGq9h7Q7poVMCVmJ+ezeo8vswrcaUYY9MHiwT7Lqu5jOtXtx9JjRo7HJPbFnK4k
1Feq5Bs0RTIV7FDtkK4SIpQicghM2hXY3dt5s9rCFQpg2D2Yysa3In2UiOT8gXIvVnZ0IjKumhJS
b6p+VQNalfA1sEKmxTcLZ4OBgkgzO7wXSbn5zFTc4AZNVGXylWmUmUclJaQMo4SIEKIzUqRXMvui
+w5u7mXcPSYKsqMrPFd968NzL2GyDEdzSQIezpEYTuO3KivF2j1kpRtFXyUX+w37g+JG6dSakqjp
16mY2CdZRA6+3A7Ak2/suHkBs+169xbi1TH7LzQCPpL/aUpK5VXg+PxOHUfdQmH1F+zbnmh1v4/N
MJPm9kxB++KSfwWdMmcvW9+dtV39ul9BCUltdfWqzFsPN3+4vBdHy3oYLQocpsR+393jRnHAh4Cv
sPezmHDvNra3WB08qW7OFeNFkmzvaHkupnm063yWt16zdcYTVoAda0sL3LCv9OpdE/HQIGIMuhgV
zirYyHNg8+NB1SiugSVmFL7AlNRULdFqUm0MAIrhNvfE/l652dPpepkUYrxD1yyXAAdA4XB2l/K9
biM+P3GXn1eDdqvT0PMbZX45d99HKVF6N7Clp3PMqzorMF8D5PlBA+GH21KiVsclgXMoANyDIRl9
/zS+FkqH9sZPyW3ygZmBqW7trhRr54j+Qw9hVxIAcEyKb1aIgWdXLnG9e3I42nyEONaBKyI/Fe2j
BPrwAdFSxx3NrvtMiS4xBKQoNo66/E+9Sm4+7c8JsVwdWsbpNl84lXUW8hj08QbwOQZuaGTxX10r
vb5Wqw/tuWPTPHSm0hWfYXM9cZ/MFfuYbcpb/c7cvbu6hA9GY0lhy1GS4wNhVyQrinxvyFpFUddB
uLBGA9Ld03a32F5CsLMwbRCfY1etVn0wmtbuovqNUYtbzksZwZ0uGxwxWa4hGXY8Gnx2cnQ/RrMT
PXpenBYJqYVv6CvXHGNbVsNznL3Ke2OnxLyQw8mVLDv+2ts9peeMbOp3yZH9SxdquqBp0oqpJeIu
UtOpXf2BM53CeyKsYdg1kBgb4N8QVCyixChrEWjN5EvJCbcphygZF/ZB2VDWMgy7OjHUBUe7qbg0
SSqdvPdmFHKC9MzAMZCWofTsuxv9F3nrWNFlD1PBatSHRJeqRSWXP5POv49k6v1CBh0GYYmmvRfE
EJ36BQMPNtlqM0BcOkdWD1iqwDXbpmOzxJNxi/NyVsiCJy/Hf1Nv1R4okyyL/LyJYjmQTv9pwe2W
XfujOxZ6jq1lUv+Q5q0uyk3cTYrpaiN8vqXak4OA/A4PqkrX/Efx8qt0CE1pzgStoHxFy47RfUI+
OKvj73OfLpobjAFtK8UwwwrygJ3H7nc9/6DJu2OjqkvyqxuuoHZXXb6UWfQ7Y22/QcQOjwyiseLm
tmJz1WvuvMLxMvWTypDocT9Xes0oB+BLPg+CW0iMaw9nf83lwXW4I2RKwjNSF4vKkCsJKVS0eQWI
1wKFlN6LBmzdMljPA+Y0hID/gx5Ikvb5V6fRu1apcKX0JKG3JCcM61ndIcsY5O8yIunFyRSxIPcV
UWtfQkaFYfqGqSntX3/dLdfcHgCoKi1hUFtOOne4KxHxJxrGDRdhS9HNzMvaNSX4DXt3olyOUOfQ
XB5dDSk8Kw4rQjfl1UGE/uhBpMtaup98G3+eQZtWG9pX4KqkrK7MuyZJYP4Pf7aZyh7udfJ0fyf9
OFQTb8FVkqDVcQosxZlXz8+TZL1+52t5Oq5DCRLxBx4h9HKxLOaOIHMG1aJ2b6m/uXog48HwJFqB
p63s7Qj2jeRYZXqA6P5zYzs5Pin/ZsO8v1dyuVJUr04OpQ3AgThBDCvdN0I+ANJcRL8SWZZsVmQZ
fv/FTgnQeQ977hqzQP6cJTGHAxiWzg7dXOCAa2hVYzNZpxQF5dzU51wonKrGfpbTaWOYZ/CmBV2S
p/zWD8Z4UINeL9zjBz8gh5I8NMCRfND/H2FG2fbe7YKrC7IoZpB1Qje4TqWLwskL4p9OwArWC/06
0Mod+i0B2lqY9t45U1Ptw3NTJRvXCdEgAN4eNDYaFJF8ANZrn+yUKQmeTwHOoj8VFsFUnlFyrxPZ
SywJuJ0Qpk8nxc560UL3v2hSqS6XD52ZKPkPhQKyEOeBGos2wAilRXJBBwCooVhxZFnAH+37xEtK
dVxvxFaglV5A4BananEX6W+7XvH5rA5i/JJDE0t7/1uvP+UeHpD/F5m+dwPdQG9gkeijqKYXnwNz
fGIcSGVgZlVKbRZRvFODqLs+cjC3mE0gtiyjxhjD04q4FmsY2NFEcIyCq2eUPcZdYDXmMSGCp7ct
vWkZVlSZ+W41p7+d35+sHMloC+7rVG2j371VOKTl6gctDkRrZDLnmr/f1wEj2A4ZdbPh4GyySFpU
snThmopLOxXpaM2pIiEWQeeikCD1qCPI0XQq2LOhagsw75xOH2b7agGYF4l7EGPByWnsz6MjpA75
lilXB9JaMsf2xDIjULL94Wyr/TvV/0lcK9NVDIFWMLKeksjhQi6sLRCSh/se4GMNbBFoAp2B7zXQ
G8aUNqm4cMwWW+vqF5hgFIHPF/oN9ZosjKRGEX4FPoXYGAHVOa9EiJVvBQlS81hQtPwIFIRJ5xzh
QX1Szusip1CQEWO4D1JbUiHc/sfZxMRBvAEKmKHzDRPNEdxsZwSCztjXlGHsuZP/T3nct5c2DAfu
oiLkiYuQE+jhCu8RPgTpiZHpNicELKRU7v/1HIXWsWzAN69pGTEvi2uAg4iEejnXSyHwj6Dx0E/a
fIdn1HyCmUKQwhDWqF0XudAr0qF/Y8AKsi70Oxg9Nh5CYMhDzLTr/Gxu9WDIx29NxnrQkVyejlFW
X81vMfzB37cRjdET6TTRFzPh5/HWO30/RHNu98wmQim2tvVTRogHCzw+3QeorWmXoM89wjHsY9va
PxX/WEe+rELy7ji6dU8dRvnx7ipSrj5XQl8NUV2G2SVRgmL3afMp8+cPjwITgIy8FCc2R3ccBQXX
a5UpUby5HVfbvxZh4fyEFW6mjL8NL5nRk412pfCXkMaJi/rU/nu8N3bWcDEiXn1eRUigLxR3z8jy
A2NXrPnHgmnv0w9PBLpLN+61yJhjeuCPYd1bjoldAFMd7OW4Wa3mTY65yZtyTJRVRIHgOLIWCFWw
ofUKy092RN7e0DggMtEbL4kwqh6n2KqQfRCBN0wSDdKsd0XfeO2duBgi//ekYG4X5T63OIbveu1b
z1MHsMWo3Qu2uYLz4863PHly4WVTrXuavBZ6ayDDz6Ws+YdmiXf0kaLopsf5qWZxxEiyfwy6ch2y
7q6Yf3ZOqSd5NI0NE4NHKFpLrZf4o9VtGQ9Ks/rxz/57IfDBRbWCI91rjN6R+XKCMnNVpESQzohi
A2iwf5HhbPP5y3pwD8he5bMKr6oqxFPBwvMKm7afFO6wP+TFS63qQo8KXrtt3vvRGtLHqyRI1JSu
RpCyyUQv0DAWybV/kKH67e4SyZbnxYLDhCqTDWpXp1okEDJhfe1/VWGPnjP0peX2JeB0SrYEHMIk
JzpOdcMAEusblY3VTdrXhZPWtz5O9GMcT/TFFNCSlhug377k+lNoMWR9CB0/GgrsZ/A3dEMk7SBI
XUFEEo+e0OGe2cXkTvILWuFrLyh1R7sXbpoDx56gjufbAhq3bfH8X/qr6Qi6Tg6jS/zR5vaRmc4H
tjsKYl0i6aTfHm7V6BXFXxqlQMEAwAhc0jicOKHGS5jMe6oNpvMaMBgKYo9gA7Gs1vk56loZqf0o
VoCeaV/6TJR3QJ6tCeVyf835kV793PB0kVv80nz72Y3qpCN3Kyn9gEHzpRmHMumegzHwNmCJUbXM
J9RWqa2V0pAy2gVmyonzFlDIHlu3hr9lSDFmwpoeFzr0BnY4F36lH1zNEZ4kjDBkheQobar2r8GI
r6yYJHi29LjD4OiON5UabvQ4E0Ajo5S4yn3yce+O/s2SP6vqGT+0gMSFKq7WfPdGNeanrvPVycqU
Dd7jFMNMXkGznCvE8GiolMOq9GUgBnYsq60l/zaGqKijgJeEZ1nO11UrSeo4YcKb5s41/MW+BoO3
qrkPQB7dTzasEgMbeI0b61GtLX05RieOoF2UkTM88kR0QZQr/08QPCU/jUgZmIITEgF32Krzalkp
VtrPOYaYNq48TX8t30n2jg/NwRkYml5acK9gFWAeKUoV9FpvXsXi/7rhwlLSZkSZdrAVyJFpIIR8
0t5pzNXwrZiWJYC248zjImWdOIP/YP2vHa+hT7XOr4CBpmTQ/ViuWg7ccw82bay1SOcNP31t+tYX
xyKKlyIncR9ZldETZsq2zlO27yoYg3bP5inzQwx3sUKV/yFWACtX4esXNojJthLnuw/cu0qstw2Y
J0islW+QkfI3vG48w/vqiEEgmXmos+q0oWeO0BRfkDgrC0bb0QgFjz7YFhstCo86rjkUcgjL7PJs
tIw/xhhGTLkb/FvHPINnwoO3Br9swCqxd0a2a/r6LYbl0Bjet59SUwfRUMnnjEDvSFVs400+reJJ
hYScvIVyEX8e5VEUf2InlrveYhuVN6Yehjy3FZePsdEM9xuQkuBc4wemo0w1NlN8I3XoSzUokV7U
rfs02i68Q9+eRdcctkTlhs9YY/72KCE3fe3ojMgVClsdCqwYF8NAiN2YwQWzH+AXaI83K+kPu9kn
+cNw4yNkPN0v0Wqy25N4qUEjOWUydy7mCl9HhHawYJtSNhec1bNwf4S1IRWisf0AUTYPJlFMGeGl
b5EzV098wu2wJuXIhqzuG4745x/ldQ0nUrFGyfBEXzHXoA5aHPsaq/lCi4JByO5a6Q9sC6vAYWfE
fceR7SdKby5hHVSHr8+RBH2HTZ00zbhXq0YMoa+GDzQKq1aeTdVfABUs/yUqGa1UKtJxZZmBQbSP
JT7f8VSN/3D9j7C8DuEEcl6DevIS65qj+qtzxhTCvfYEq51+x13y1birX6iRdlcVlutR1oVlwFG1
pYlRXdC0cVGK/mo7J+fsbr+P7DTYawUVPjegXR7Rp6bNK9ZqtniuwXzC8F1xoshBnM6g6X+7mOQh
EVyiVZppGil26J993aVMucdDVamoh9CrrGQS/rdZm09vot9j71+NaZ+AOp/zk94ZWzSMxJ6IsIc0
hsXz8wokhSaSOBZzaWTUwKqBo7u8MprDIYFt0rrfo9nGdccsg03474CEo0/BxLvhqeCzD7kYahxj
0rK26wrEfJmRTvBpQojQ1CtfT6WrsWDES/ZjQIu4i5T00u9f0At3GVS8SeVc1eIpuepXPPj3b9FB
QF5EXArtyvawbVYzfdxUdZfXw1W6BF4LP2r105N7/hMDQkbWQ6s7VHjd3oi3JmJVJBwdS0X/+HLp
b/I4+g96MnJHZd/9yKI7u5vvd3OWKTfclhUeoflhbxsi76kTqH91UKflC5NNqIvo4fs4+1ZT9qBr
pxIRrb01MzTsMB9MbWeB8fOBsXnl5RhmXAwHmEH3MBxkigob0qEHrFFDp3Omc3AO96mUcm//DybC
iZw0K2uAAu1KV37oNMZ0D+ojQQ61auEAe3xiJZBrRXXHwNqkChF7zRo1emSsNIM9iAY/VtNon8CT
aO+FxoiCELkO4dzhDIZAbhxyj3CqL3SX2gBVe2FL+zUIxxJ4fNFQ1oAIp6m1f7eMKnniI9PtYazv
jFZAeuDjrvcSRBTNfQzb5oQmhOtpwwiAlSHp1QO+7mjiN405IbKoEh1a7THC4O8yLsNrhjbi7xbY
kr0Ef5Ha/R1Bw/EuJqRcrjhfKmdg0FYozOGcDx34buKBEK7TqM9Qt2+0Uqte7xQWavSsRQnlsYZ6
7mS3GqFys9W/ALAPCapCiZRhzLbXbLFlytIQxK610x8t/CVrhU2HbzZlu8B8HaXzgeOEQJolTlFO
lQELiyiwQGzzmzg+ZjU/zhL5/Tj5prTiXHB4QSK0bCIj32EQKP70KrOYXIqVl+jfOuUBkBcVXxbF
C+Z/GGHlaFQbJqfYQKQmv6H8XqxhbBG8M+oP95RwlO6FV/aquW+Xum/4OHss5lJELMaQRfIVFBro
hFbKRDevuWC1avICT2oCBeO9b/3JS2u29BFT1HaGSlrCowEnu4Juo3K82vWU2ZDQSoGhMFDeAlqq
x8AfhcTwczeK0caqLHrc5WPh8y2Z9OybMJ+2NmQ3ry6FwJUIV2wru7njuGFMKjVbyqzx4m2k6Pgz
Gijb8ZDBnRqOU/Q19xe3XahTmcfZ1OUlFMRVftXravNhsDIKS2E/IKn94OKSgi1wS8PoDUr/W9yL
WiD/vjL1je1EgoWz2C2y0F+d9eF5z59MDx8Jjo3GlNhd5vWhBHC3BIcS7hcEuiMYr1dsVXfstX+S
q9XeGrh5PGb7lhzddzualml85LKUv20/b77zWrZLdn9ZiCnZT1THKl2KhJpl6mhk6Z6nO8ESaoTa
CifgLPpZtW7ApNQhYcAJdLca2Cs4pmcCYPbK09JQjctH7k5ULOdq8Nvv8SOypXQ89FMT+TfY4sTq
aF/+HdZiF1S7AZHiDA1CxKiaaJvc2+DS1AsZNgj6OKlg0VNhUVeFN67xn2kpsNDHMTUyWFW9mCYL
5q8WTyBghIT3Rs9pWwfopZQ/N63cfGKdxx/IWxgkXWqdegiAyLMgqrPtxqVOBXm3LkKEyolGQwKO
Ulw0TzTcrx2pnTTuDLbdpYFzMSpP+V6H7DAcslZb7YJxbjLCQ/cyCCUq5E2DY0G5eUy+4Jne82kW
fYxo3UsimonnqKSsjHlNcEmWqAqlYPbcMb+jGfTqpO6PtlisQiVG+FXTx1ahEWT6fAE6HbsuVahh
UGxIiHMrCHfH2RmNx246Cvgq+bB0pLvC0SmaeTtJ2ozOUbCQB1rwDvLTLZTIKy4JtN0SxXxT2y6S
GR+WeubSRclGPG8cGRi/hoXM1VOYy7FhUAU/nWvZtDishOGID0z38hvPGPAbvD9kwjAVbQSAACDv
0DV/SyMoW7VcavtPl6NumDDGyii69qiUqGBFkWT+Q6R26MonCP6pufdnpI+C0uxX/3CT2Lvm4qBz
EUnf/o7lEMOOjl1Vc/p37shDS3aPkH4gziLE+fF003GxJEqaQWflFTJNFYG6d0l978tJvozUpK38
E/bpY+BJSkT+UlVGCTIKLdRbv0OSlRYtpfbfEb9JCShMfxneq2JRD2VqWpxx8l5Xpm6cCAJP0rsE
6tgDu8wW4RuqdEii5pTLFoGXq0XAhgxIj7FsVt1e1wxCRdtI/mM8tTfB4mbBucicwXdM7Wm1fqj1
XR6f/JbCyshmBB5hCl7xdmye04wYMOQsKUG0Yby80ltIcuTsQ6W9A6eHCy4Lgif2ewD6NTb41E1j
c7qAlMQ/qylKWYzSDepMFYQEn65A1FUUbTt8gyQUbSBg2pbEsddov5HpFoxxjju4J3Qw1cazH3qV
vY+BNGBvaroqfxAVMdvHKGjCeFN/evfz4tH0MBO0X9YmAEvZYImV+A3jPUzuoKYEIw/vjK5yzTua
JD+2RVrKz2jjxMM0WFOlnjCdsdEsJG/pp2ctCmyIECTg8ZXY2GawVzG8CBUPjqLCkAlom1xKPyXC
sfAG55YeTlH00u1mYoT1yzOME3Cb2ru+CN3cXQWjCMFSdHoG5gPmDBWLcBs25xa1d3Sy/avcHWct
G/ItZLJJKV8FTe38W/j7nY4nqBBrpmypxmdCxFJr0NHdjRIfiaYCQkacQYEtahJjwJXaFj30b3Ow
28PmRIqNGE8z2aibrLtMI2zQQeGiL8egocI1Y4WvolCYCNcK1RadTKGQhiNUEXN+b2pYwh+yz63s
cMv9bxVGyt3UtHoqRmJtOxGIpUFI+11UJWyuRPoP+ycA2mimnShHE6WzN7/VWx/GSygacCsp3utP
05vxQsAuG+vDqn0XNOnJjeqCabeaa5hixZeqZZss2y2rSqNS1SSdOFZ3ruvHm2wjQ69vkvz2QSbN
JaOj8U8UX2n6kV2ITnqfljn7ASVVpDMCUFNIcirbyHPbklJeoLS511S2EuwUY94uH/QjhjEsTEys
PSdiA79I8DNCXsqh/ZFd8L8HYx0WFfFucjgVWIjZyg4z1bZwYPHJ1OUv3k07+lLO/1gVfWyaUvVR
uUldBehIpcw0/D7ICZZoj23s0OF6lOSBCoXCtrixguaaFlDkIYF13rDxWH4xyfQwlcocK7d+jefS
bNNmytIYSn3oCNNoZLG5Qr5f0qiz41EpI1Vc/zjBlsRM7/u5cmCBEdNHkOZgcYO4Hye2QLPIXCj8
m6I12g3YU0wsbgL2VV9dwWctVuLwjf2i20Vfil3p8WCO5yGTHioO9DxZ8lXs0+qkignru2rbIs24
8JK9q2+w+qOXDz/dBSGh01FYHon8mCn2wumDRjejA/1ws5T5+BJxzVZdt24lPo2ICbi8G0g+l1j1
sbNoCV2UexKXAp0m9Eg4YY3b74xhjG8G0Z/RUFr6xViAN6S4C1olPh9/iJOXcVE5oijWjemLdzYT
pbmdW/TU5Dx4nX15GyX36xoSD9/dQXmDG9IQ2lZ4+T+at4ftiI9H0Kui4O3Kve7IhaKhS/mKzNHs
oCPkIgv15qgHu+eedAmIqPIxekFlIBqER+IY+abb5uoagqNi408/7I5i+yktUqQc4mwe3ILS4N4T
J+m0nVY6o+hb8BUdrjPQ49/iDZNxKuEf0DnvqYS7F8gL5LJbtlZ2wieDEaTKVFHdHBfp3xMeQMyv
d8U6uNTxhkgNLjtA0ZTX0fFfMdn9wVHpynmGbLH6rtyIRWrV/rcnULiFxA+NgylXraZO5eVEY/Dg
Hu7uiPKNZKf483KQEukN78BsdjANIVhG0GOn9H1l47eDIaAhri+0hNaLuJGw5UKeNxvVNYwbOJn9
OFJEzLE2A0O5uDuCRPVDZ6TlAbiXVASOMip8kOsJVkVqlNCAzq8T24LLHhLzFukC090AzpDZohvq
H0a2c7QK4DByauBdTpFYlhDQG4CjYSrUESM9Gk8mT90k7/8mLtGIvwXvMkWaDEMGTjen5EG9F9eZ
9aTzGVsaKBmRwr8VSzFBCDUxmSdTWWlJLY0zvHWAh+EcXjjixJrsUO5WNCCcKAEeyRfOj1GaO9En
Wt2PW9mosfUQfa+W24COfmblElxWB16uXbzV3bQb+buvMlSJrB7tYU0/QJA+pWg5Yqvpc+v+Xt42
CIpIAYNYyzk8Yq5WzbEyiVfPNqI6eJXwT/VAdz0qdkqHqBV9WAZTbXAth0ln1wmF4BlK+tyAV4yl
V+LkAY99ydfQCFgYPNJ/nrB9Hpd7YvNB5qcMXjeZoI91B3y7Q8mJunXcEgphnbXg0X3GiZ1n9Clw
oqedoygoORMcZLk11hXpXzT7xe2kTSH7iPYqb/LBBoX7j8ZbF4Kk8yIxxjSUx9Xl/Y0TSONpdF52
qg9dLCD4T0vK3cATZxvpBQUGPi6pX063EYayjGPSBvzGpGlBW1VfvwlB0ELVX8mQHxtVndkvAPOA
DXBlUWtpeD2+F4ZVLWQICicy6o8OMjmjrc9y0dZuG6XRpaI4Z9rfAB6y3hyPXvW6OU9NAG69mTJq
VcW9Xs963f1LuxofoRlAf/qtBfH0oCLUw7y2hIpt2cM5Jl9YjzCeoNN2Tg8LClQEVYerw3dLdHZW
DU2Zwa4R1r0iJNaq46Qmor06OJ/O87cUna13UhQ97xfwGrWD1WZO3C+Dhod5KpIN1vO9MZ9TNWQ9
SlNHm0aI4b6UBvOsQ6obmbUY4JfNhsspcHnJTHG4T6eu70vv7q9m7LUdgUKtY/U008opz5uakodB
tPPXfoKihll2IcwnBj+V7Qatn6pyBxW6PInOX32lytSal1BNcqf0tq1Y5OdGtNwbAbuhRQ2jsav1
QTHGCx+h9DjbN3w+TQN8nbRXb/8tKXw2+Opfaujsi1EaheECmhEwR1Zvk+e/trx26LKb6hUKc726
iA7Xq5l+2q47u+39lFotTrUAda2McmjwzwKZwyzv+trPLw1MUqzfWAavmMH99oSILUs+WEuBuGrX
utug1CEgYPZUrbevgBRNRnmvJHaT7QkSLotJa9Z+OtypXAS9iF3pLa2kfV8WGd+Nzz0TZSipFEZO
DFcoYAON/CX4Fj88Qx7/F0kTLxBOc7bWH0Q4JbSjqOmPgz7baxt5nzS3pKk+qbkhXO7wyyBEIy8u
49FYWtEA3wC14x1TsQICY7H91rWGla2VFIOaj9DIZh36KvXGTs1Ue6LM399Ztw2fVtdrkYSoc/yj
0N3PJOoMShYiJRixhS7gvAH5/lJU0/vP7/BinSrws3HOB/00DzsJhIJIaGV5OTrA523zP7D7I3ss
C7TnGpcV1yThn5BVi3KVTB9Huf+VgoeBuKCq2akAJXCcobcHT5WAvUmRX0hMBql0kUBHszx9O0oG
UK8g4JeKpGLp8mnDSGuVjQBrCWL7Jfsm300X4SqWrUexal/xGQw1E/7RBNipDxIJyRNJfnNaO8DT
SsQ/bYiHVIH6YAf0zZ8V7ftAupACDrjwBwVh4MaIUIMQ7lHGEt/BNsPrdHFmxcDq0xeJhtUjcnbW
GvklEGh/zFjh4FqhRw2c1KGQk/FzjSPh/nk+HsGNj62DVqVP1eay2WtofAt6BJsW/rf0+oNqmdHS
tbd12cKNN0FY4SZrUTCI9uyMyMlByAq9tCp61GnXYOJUN+aGa2kKRRTOMX0Ogx5bh65En6UAD7Sl
OOjnHsmHw2cArJqbZJU5zAScLseKFi4Jfu45e0Fu+ensl38vEafD93/k86oO+QL2tm4YK+FaN1tA
D9hnKJfGWI22RSNTnOgkSumIW6KvKv66HcTDRkTCDsnrSiCPvlhb+WPtL7oHEfOxaTo4nRr0h5R/
deiPOxR7/W9BRWfj/xbr+xgczbPhb+qSELLyPgFOu/GLe2p2Jkqrkjb3kjhfVCfPbLA9qHE1oRAB
/mV86HRWd48q0lKNzm9tADsANxKd85jFjB+fM9g8lP/llV6cfC7/RMVHKon6tdhCz/vis9h7VUKx
WiqTNQd2wtU5Tttnid5yibZfaWhhBRoaeTz+ffnJw1axKqjsaggIIvfKxQK28ptKUBCF9NM4yNPH
s8a23VJ5uqh/ZHR9fGbTu4XwDMpHSQF+UVPbYNUkGbQBZR3YYopj4r7IgTkJrJUNLwZ+1E/HslE5
gePyATtHT6ggFwetcLXOqZWLuPtFq4mvoheD9o9IBV6kS/7XJdUd/X128LKGY4zzjW+V5CmSvpL/
dCKqu5VHspQAJZiaBW0PEBskZFGVXZqDGwDwUbStBU1jBzv0TLDkMc9XJqhB7JTu6+EEmDJM9D2i
iqWfHkF1Xnrro/bBoccMUvj9+t40C6anr1IOmlI1qJVB+Ub3q1oG+aR7UTlwv1nIpJriXjLk5dqS
6uX6cJEvNz3ZrX7dRbtnI7nG5W8EweVTS93tsT/TvhHhmxLKVPNhA2HnRvoWGbJGwsfTia8sdLUf
IuO1LH4Ciz0T7jS2fxqyGCwVxjCbytsfYKwYCQa47qfHyzqiPTKjz2Qh9fGqYXj/MxoXAzMXz4nb
Q0qRjidkbjoOfj/kaT0ul3WmTwdpSTrxXbxudZfcvN/humugWQowTU56lchbeZHegP4iI2dORECW
/ONgt1if4XdFoi8sielnNG6s8b4zxO21Rs/Mr1OCBNlkfrboluE+lXRPcFxmEyiUa3BuVZBNuuRq
LyTHPoZCueXmaqCx5V5pIp12lY5sOKzg0by1RCYIxMk7YbLrm3l6WbgIozTNt7xKB/NKa2ChJhub
LBcnCVdIies+phWHvIa5quvcp9VA6QBmaHdTXESyBrBO/qbV7UrzkBM8umuQshnaQnpsfA8xbayV
IyhlBvg2v+BwNNHyEB6t2tTB0Z1Z4Uu5CGoCu5eE2vgMAwpwou+9fAwkTtTklcvSfXo0N2JbwajA
1LYmRdDlnt96zln4uPBKOEIzbPS5cOjI3aoU2ErLAMxydQYR79LARwXlXu1DGkb9A9fVR2T6b6eJ
x35BIXSDIbNoHGJEH1b+ew2UzTau/ZqymLsVMw9LWR/40mT9iyNbOBiw52iZBIgyIk6k+woJE5qj
9+hBREfXbBeF+jy3c5ima6oPScZzvfDomGoHx/znozwgcL4QOHZw7WfbytPp6OxC6gfcmXf+QxlK
cWIx5NVJl+dvNB3MFQVgYTItTVdfqBYa72bsHmWEexattRKkRcCOZ8x3WjdxJxBIH3kb97pAiiZf
coUZU48pw4n0uQS0BnUvcW7s8e/c8UVeFeYmmXpg9CBS3TtYrBvoj1JnG/1m8yn+NE44ykXZ567B
lHfRfwG4iEST/36fu6XmsJiqJPMhowdshbnEjtfwTNGY2vJQzDBPTkBcBNLn8zfHv33jmwPhHEfR
2ZiFH3Q9E5WcR3bLW/KAslEdiXvdl1h4u02H/a8dGKOhBsHFxP3Y0ORxceExwMWxBYL2ZiPCQi0Z
wKdwkSNiLPrZeIM8YQVeKWzVmoSujQp0ZiATtsCGr+woLLC1wGgXGVYt4Jtj51+0Bh3vrFErnupJ
tlT8OlBcq2KAKdKSn8bNwLfp/10YOenadJHFFCzQXd1tRjfHvGYcuAOWhz1rZptJgDXq8aAIIpKK
9mPwA+N9+5360eW3zCJY4jRU3EJ//PfQB5p6zbgYt+e+GHzWx+niZZidoobfm2OJ3F5S8mSfoZyX
hjm3SPlKSeXQG7Eq8qtusWdvbHBhdgfG0PySJ91IZRC0LtiulC4h+afR8U2VH1KW2FnwBvHJGWF1
aSNtWQHMtpfFYGs491s91ZyCNOXG6zTSohCeRiI9cegw1564+hY4gfE7fkymjN1dSkviHyNanhb0
02080tOouMki/UI0thUBESVuSRUo3vVLXq6FXsuDVMRLkoxoEAhUB+xRfOyWZkhXVpLIyLMwvn7J
3hfs5sqeNqtafpuTAcQoYUP6N/EZZp/THjuwzb2ThAFmnB4w0Q9RU0tsnnjaXdZiASLvitbO9Vwg
QmzEW/joGVfXlzDJk/hTz3KFqMEKzTREzT42MTxHHvN/AGurJ7vJVTcpUfoyFMcoKVYoFYBY18Vi
obtTySAsuS+YMSx+bRg2aYeyi6l67IB2MI4EJ8KvYtWCxrGyVapS1I+pEfSOoKj1OBtJh4Xp3pVB
br4dv1YcvkPOqPoC56TYVMmUeRljWb9XOyQx9UXnR8hvCQ4nGUN6FaNEMRnJuIwn9uH8qz4W5uGY
+2+4YAFl9KEBbZLl9ZwzNHkGDqCzD+XZH98kPtJ3k9kEMG5P9mkjeuwsF7hnOz7cuI00SKOyepz4
wy3fzYOSts93i7vTP+E3w1BLau57yr7UB9nR1Rhvwpzcm1UUzoiRPO5IHEh19SGou7r4H5e4iJl4
C5U2OenQl8e3fhcPLmjWi2Bjsc7skkr81oIHZF06Wi4SoZVJw662nxhJ+4ZweSi0rmY/kSX1Lhz3
1XbzYIIybK/GHdov/wgNMgNKVbqsrfihw3MQ/+Z+OO6LiWEsfCJ2te4IfRsPUULqU/oWbC5wEAI1
EHCXidPx3LgukxW2JnZ4DzxveLpuT7QY9AybwyIgIr69dsBD56c8Nqbn3iHf/qgUTUX6RICcIzMw
Yr3sU2/T0rL+QG2TnygO6faa0zxhgnV78oRh+hJBeJsRviMwRmeFgHC/1Urlcb1/713U6UDnhzCm
19EhkDvVTj8r/U7rED2JaxSpTBgsybiaxd6NWyHzkvSfkiWWtGziImvhabqEOWO0LdoC4+Z7Fq9Z
BnMmTcNSkw/iQtXbcoKfZTWEeo5CNZ+G5sKFk81Hpmm9nR69LpisS6gZwFt8nidAe7GHiInV6ocZ
g8sPH93wCUwV0TbD3z3zkOOStOcP3zJ6GN7dpVz/XzLNqam00n06C7FBgWGw9yE1Mc+UzWkjZ6V9
GwbOqpKm9g0jXN6Oi5GyZCpwwi27n76juVolOcYf7toTpuyTWDXEyeQ7OAFc4VmoLW3Bpmf/DNR5
lM42oxRGxMbjtKfHAVIOVQJB2vCC67xaitK+eh5/t0JoUiHuIdF2X/uxAdMtckRdz4wCsFm183q+
4HSjlmh+sqDyrGSrlD1edxfeFtGtM0yjFv8mDlo953SKttLtlR2rgPLTtjDzmO+M07fpg9B641Sq
0CrTDfZIjcXSiiEeS2e6SZbQCetVcsAI0S7xhq2iA5TJ63162mf2amOwE3QumQJFFz4kuzmW+1C6
TP9/j0M3M18cWrMJGSnK3ku3aRgImPYycGqM7NEjhg+mTGbF/eHO062GYqeYjkC8iceRHNjf/Vin
jZm+A+C10QDafDw+04rfgIOSBgl1c3WcAXLqMsbTznD06nLp57ZSzdqqYxFP0gF55bbmLrlr8KBD
nB3SX7caEdKt1u81fmbelHprIhHU4XZ5ZrfTvgB5LcqY0X49FUMm3vDZFdefkWXTifbGFCKN2Bl7
XTycawhreX8UliBji2rZogCScrqjZv+Yim/YgQv+r+0Y8BWYZrgMvsIBklpebR5tLoe+kvQeGSGm
Fq5QIKP2L0Zh1awHRmBveTmXOBLUiCVg/SaGd8sZliGqOAP9NK/NnCie2F0DO491SIeXUpVizhPw
YSp6/ui04GxI4ht/GOuMxEwbHo2uLJvZ3ZMdniaGzN3XARkTEVI7BXl3h8ampH7Wx4H5qS8Gczjy
1ZoTVFF90lsXddJfO6npiXjB/K3WZG74sakAyb/3KZ6PpYuiciOvNqVvY+k9nojPsl3CQQ5EhjMe
iNBW2QNArVlq5JgJg1f8ciYSKc7a91gMxebgT5SkQI9+NY1YE/sl62GfJZ1m8W68ZxAWg4xf0217
lvSQeTvyWNG5Xk9mFh3ZEYV5o+Ac6+Qcndv9LXesqq+BSkzCO+OoqJ3W5VsovNOXyRBDCjvBYAeP
RorGPZBEipyVEVyjAtWwkGC5+/dYxng4BBI8lM2jWdMjt3aK8FMhQpex9yLQ7+fK2dCGqkgULhbm
juXsf5zyP1x47dx3wdmykRjLdmgAUh3leWCE66HaLnETDd92+IdCi3sQRwuuC0Y/9H//Vt95pCzy
uYMbyvUHkAOixke/yENblWnqYgojkrzABvxaMWXHoQgcywpZLIBvjSeKXUZT974v6icdIh/99It6
tt/ZDDxl1Hp6PbJ5zHTpG2RJguPdojBUkasdLhKBeaPFTv3vNlmzagiXw16XYo5deKg8YD2zjxjQ
PI+m4pIIju+ZMzxWGSPPGq2Mc4BJ95mD6z8bnNR2tObq3vlERRBkjcaGyQ6ArjlktvWaDu5G3qnL
C6TIEApUfkRUXZVELh81qaVrLOmEfsMtfSFEVriyF6k0lmzErc8PzKiR1oL1m4N2OL5sXjdX8dk4
LM0031/URMixJDNQdefaWJKkeLTr7/rWj9H62PUjN1SlVjg0aB63UA8x8IigGGJ2vcoq7H/lyZQV
Q9e03Yo7fd1BsOU6ExN+Dzd5z2q+iHtYIDYPShTuJFM1mw/ZXyn9nRBXhJoPUxnxwo49WvSlI8lu
ZR/7Dj0bZao80Yg88a5y10GkWgjUtLNlB+BUnr5raPpbj3HUqR+JsBTfoLrx1K6r86ANXoCGjNtq
NtoCWAFs7+i3+b62L0SOXWbBCpOmrUQXivllWU5VLZg9M3nPzDNW6XwuqigsWq03mUGmhty53O3Y
7FfO/xmCgjQhjQ9a1P625bw2+RWi0Fb0HbPEPGYTTYoKYf01FatL/RJvHFvTsA8y8YIKlTE1ohDr
HYa/yMq/FHQMFDY9v+UaFJ+oF4Y9tERI6rkUaFiFODeh7/StTkBmswIYy9f3BDWuDCWjT0j6M3CV
7yhfM/fzpdw0oLaKCPTI/iOAhUDidx4PEfds92rcR8NfHD/drGY5kh/cnPfPFg572lco+JcMvtnS
w67LMdtnJeT2gw93xRd4/liw8zF1Q3pA/W32uTEO1eXkCPXYJGdYgJRlUIaJFjLYa89jiXmw4U3x
hzbrnPZ2ViEr2Rxv9gcD26GyMGq0pbrioFfekIH2aWBZJOvi8JrGWBdOUIVDKxtWdoWgU53PkM/j
KDxhISk9/XitOha+MEwTZFi+pAfugKte53qaxoQgolpPLv2947JNOXmvAhFoRnnwHtFe5rTOphVL
KNUs1nqc5Gptweb4yKSp5OVsLclXtEqmVmfCpUXWpcnuxLIzIgSn/T997fh3t6xesW+srmU+AWmM
m2ln606Oe4MGsZnRUBlogkEBMc3SlPd3szstzZSHxVN+u6pNofoxNZ02o4m2N8OKLHNFMAgIJqTB
CuVumr7NBZH7QD/WsnxmPWrRBZ2QoyAAzXrCPjcZxg5Q8YbKofdTtNTWXGFyAObmX22//y6cU8SZ
TgG3Fyd64ItqSi5aM97XC+jkXp81wpQ3EnJuqoUUDE1Uw3LpsRHUyCa4W0XHFrjdCU/GbDfPLT7D
+Vy13T1ZK3VAkNuErx7TruxZpH5OsUyMhHAEVsBKsBUDidBGOI4wTTpS09wCLdTPBrQRnP9wNZxL
Lx4Ro4huoAar0cpq3tlCa8RdToJJG/ljlHrJwG+J2q3eRR71sAsW/vDwsnl3drKw3w0v7xSzg50E
F+rKjAUbTx9eYpcsd7yObyPEWH9MsFMHLVci2wkLESX809mL3EKcPOacKda+GJlYo5ja5h6YxP0L
bja3RR6f72SE+FhHVtlZUjLZKHJ/uuOQ0kyNZpMp1QhGebwDlyzQO9rjjfteB936HWrU5J44vzXr
v3Z6KNpp7NajBVVVZ4xVgaeuwy80ffbc4vMgKe2eLvCls8g4jNAzaGLjJfbcRl8E4cEMyZLFgYK5
NqFP65Cqvph9/plTlHxp+CqOog0GBTddf57d6FMdI9MBGqh3o7Dc6GNvAIHJNyB1v/WraGXTTgsD
XKmoyMV+LhptXXIVIJtc2WTetJSVqaVP/3fl7S9noDcyId7+XH0tx/CIXsiGtxTHqymuWP/fA/uz
hr9uMImXsTn/tTF46uYshlLJ29PVoBbE5BGi6Ku9jcmiWmbORs3tR8vLYXqhy/6AbxMYgWwDMhZw
nUBP2Gp1GOV5iraA8WJ0KH3eJGnJ2p/HqpiHBoXONG/JDEI+sQ6BcoG1ES6w8rLWuAc7rfFmEzUg
g5qEiiwso69VQd74/zpAn97NIN3VGK/rGAzFxz+el+r/3vlHGynaRirKUFMU2q1Z8ZjAit64TDHD
qUMX0K+zsqsm9aP/nZ4QtarIGiTD9NbH2YNjKP2XSbhHdUruvpppYtgr3DnDvO1oq7psrTaQm0Sv
Nyaa1WbPWgztX82m3Fs9VX41Rq/EydBZ4ciYBFyhGSVjxk3aBi6Go9nVMz8A6tiO0uYvdqNYrM+b
nniqwiOOjbgG4iFYGHNd7bt7zYkGuQzDaR6SlC3EnRnmKlFfdjNWc/M1W6vp+RB24kl7nco+ZQo5
ilzwZeUbWIRPRrReCOqvpzRBpvwnBB46x5KvYCJ+yyqp43s5OT/In54t05FZolw59NoE6bt40G2d
9zx9uVrz0crsSLw3YJp39CTmUV83qHgOpRjSDXXWaPesxXNVlpdgCy4OiCRsHcXsoIP9qNUcXr4l
XEEk+gbGuf9L3/FBOvFt5zHMBjGEAH3esxbEIK1EGLDckVRppoyC+rgepN/5Hh3j5al24TxEEBXH
vcXCLeTTyqgyaymwhTVEejUFZG2c2jxHHCLyHl0GjbyHfIpTJpSdof5EA1UgWH0FgmPSjWxbALj9
YPyxG1P0YDcsp3C83ksL1JWzFoQtdN7lPbgyvRdBeOgOenTxCltqRZOcDy6DBpF3FhSFeq9faBzG
gyLOt8eMtbiCeGlr3On7gbuqe7K/7V0qhWuSj6COegFSi+B4pZ3SHP3kYjdJXIfc3ub7rF8ZxEYH
5wiCeDHtJB6luaxFMyLXWUdaZLLWeUCXWEOZCK1L6uBFSmaWL9IKS39AfbACzwB8a0liI2926oHS
eTiKjNUKQXb8QalNraMS/xk0SaK149B2f00UH7nQQW5Btj1FA2+GQMKKvAj0AB98kzYuLas2j4PJ
DkVgDzsVgRQ3EuGxwmo/++NELcDlwbtOhwxS4GskxZw62TbRI1VosEYUFLlM/hAgizrKuSbxQYHP
TTRNwxc0XrejulIxqi73/XSrDVu+z2gPkV7nkmtEu0T7YPr7iXGt/FdtSDiX2ZlplARcUeG7e2zY
cwfoeqWlg+uhjdc2fDP+Hul8FtMDTGwHU4SEMfnVklaMlttKjTVG0aZZtcjeu8P5sXo5slgRueGG
UnS6CmN43x0sSRgIZ+aCaPwB+6dTF/jHrAVtT4ME+8GLpgyIXohIiOmUPZhkm27WcxOtx1z3O5oO
Wp78k1z80ebK8x8t2y3tw4r37ltVWtCzV+JgICrEXHOLnjbrJHJJmkwzGAnAhpGExbCnTCViGGlr
EzG6Q5RB5aOlhxLxvvMTuuaZchVkHJHz0zdwQAOtQCOd0R68MPuVgjk30RdTxQ7imXv8CX5kMQaD
SmbGRNs5x4HqifytITfSCwWlR8c1s2PSitX2p+NW2LzxwUXnCIHSpT1KjyZ5pNFmj1Aoc6D/5TCC
Ws7Cio+W7MIU1C4uriGF9r3ukOQYKJ9vNRB0KznFdI8x/AXr4ZxWqQ5CH8eWvPFU9VdHN9Gk4HnP
sePeterN20gaqrqspByrkvHClm9M+eXqfdTAX/Ovf9TDGpHnfTV37oEUKVhMxy5/NvR0ofYmSqEJ
6BbE6rLkLvWa8EHPYGdzDzaR6/cSVQ+kK4yMde9oez3zAAHom1KtLN7HsyW/hjpU7zmRm+ViB7bd
5vFBgbem+pJ4X2Gl1n/bLE3JNHotdkL/hM0Z9QkborE89Hk5R18pke8FfyxUA/jZYgFGt1zgbH7L
nyAou5A7N2aIh09bUS2CheblLRuoOkQWgBx5cfzK1GAlFf4TnBrmkoiKZqxKiln8R2vif0hJOGxN
JuowOF+K9OjsmIpqgYPnTp0Tuw5ZCRexr8c4ZK2G5V5n7F2dZT+NmylGHIHBumUDpKQ3RhK76VYt
7hYBK1QXmkoOlpzhU/yk7XkrJ76l/m+jVoKjtYq5ZdsRzBTtFIEKAuw7AZzFeqk4F5564ueCiUew
x0MDJd5xiR7JJ/wWuP656dtADVvTH3CrZ4RREhXmrtwkiYzLMMYgD4kEuzF6KopuklmDaS3YHmvH
Dxy1L3uaXicfE3tYTxPL7N0XL4rxSp0o8o1wGf21wER7dOiz1PnFxZ5SC6f2FjmYBJ/NUoz3dixo
mqJmDO9SdhDEZTI6ktNyvoCDO5LxiPhM1qSSTcSPHxPmPT9LbcNf+yML7c1nBo2ZQ3Q2q8zx3Xg0
liiha7vutihanPhPFcY4kD6VXo4pk0UFZ+8eRIWekg15S+eLKhaizgnROo7gs/f8U1q0lQ3uZ5+y
rYiDSuXS/W7KVbcYryEga4DrP1J/QPsJzgZIX9SsMko3SQPA/K2YfSkJ3BP+KcTKH868M1FsCSPd
M7yn67HGxNm/McXe5sP1yJ9IbBIAXeY7hAecHpAMwifVHKiOJ3dCrcWcaTBEFeDBfkg2VyPe8+SZ
p1Dk7ZehDSgfhGJLQqQ2klAhF9kbWo3wldpMVzy7L9lY69m0diKnS6859Rja2ExLznHCEyp691bX
8Jle6T/GwoUY0VEb7engz6iSrW+BXr6K4xK3zH+V/mHjUT+J+6rR8R8H8WUc/3YSYz95v+YAEDJR
48zQux8FJsvq+bujs/0Diq2dLrBkeLh+P/3TNf6TfK0Qrf4pY3+xsuOiT1IWh6kRIsUV/myn7lMN
mrg0CXvehOS5WPFpomU5iXmcgJW718jbW8agHKgr+Gm/ql3toFEg83D/7Xaf6j1FSfamh/b+jO/+
eqef+uVj7wOLt2szeYxZSVKCqTTEsWYUU+M9nWsY24RAmZR4yRVpIwYfZJi8mPN0SRtxXLPLrKsD
9Amg4VTyWQbuDomjSUIfgwfS+IIIv1POb3Z+AXvAYg+eBBSHv2TLeYyJ9CBW0kriiW/L0c7LTaXm
IyEK5HceNyzb5qIQbC3MplMZzeh5CK8sCCId/wo6j4iwOUmTpKiBd7EXVXINPFORwcs9G4YCi2D6
4sGSG1Yos0Y0lH3NgQjv1iRy1rqM2HWHWhQI6a1vX0d4YBD9iS1MtKD4TomUEwct3I1/rit+fcKM
SwliEY1Vb9oLqpyP296Fvl9ZmkKtDKOE/QGYpX8XOmfGlWRr/0UvGgxSSjIhHk24GhbTaAGJkgLm
83qfFEbRQvxNc2p+gdCDCO+TU5aXwMjjSiGmHPugzPfQgtJJpTYLo/k0OFzbql8tuZ2Zyo9WgbV5
a2yx6wh3Mm6f3MnHSozOzeTb1vu6SfXjLyT6IkKu/psdl/DSQqdnlevgDwcUYjELewJ1KhbjB+t+
aFZz9A6Loe9X9WI1lj6SX6UrszoIQub5WVVqsVDaP75eK21aPdd5z5LXq71knsfJrtMM9dW6QquG
Lgwdi703Z2zHJ+gVTmhAcS86il9fl0cUVnBNPfA64CbRKiWlt1jahGZPlDowWe4b47cOGWvIYIve
AiHffGthk3fVVUfXsEOIYK0SEFlDu9QLbSrAggXgbex2W8YvvfTzDYpjQUCPh27/kNDTRQiloRo5
/1kCfTuGe+XlSiIfANQrgaSs4GX6UnTo+OGLRzpMOWJt83FZDePYh3pyiHvLq7nuBZJ85lKu/M7I
/Abtbw2TPIvpA3fA/7EltDmVuXgF82fwvaHOFoNZa26UkthluNC+omhxQXX19lAZVxszGkjrXT5m
24BP//Gv+ENyhm0E8hsT9uQUgry6VnLrcafllWFnJ7HDxMgR2o3RckjFOqdaxL+4bNryXisVGa5r
o5/U0ql3ZuF8EdFTJhgWimDKm5gUvtMQaAo1pDCsFrHzcLWueZtUFhHTeysiwe5QQGbOGCoYOWnx
B21BOReIGsVZHnWiIWUc935AGRunZsuYVOUBNFTXBj23My5uxcuen3qRsiyyZJ5d6AHHu/FumHyQ
75XnlwHwu0N/2trv+ETJODbkZScPhYj+hzrc4Hy+3H+Z2kjnDLbHKwGYSFUr32QCwhUwQ5fwr7tk
eoh2xCEKMg7sk+O/SQ98+Lg8NxyNOrIUOlkdOJKxjcoj+3TvsXcFmfTe+fZ6RfX5JYL0sjxaOxqv
PcQFZi1skaJHsV8dRRVJ/yL50+LX1+jjbALw7Xhe2JKfGTU3e4zTmobDJPPAuVX6B9g9r+OQK0PK
/fyf/GQhXE9Es5EKbgBzBTeRic3x87Ls6geCEViZfrv6DPVTKbvtw7A/TzqUEanGCoTMafes7XgM
HgPdppf9H/S7OKKHJ7mA/kkbyHe54X0Wjt6PAIWgtf5d+Unsr65hh15V9SJ2mjN1ShYVrSH+mZJ9
UnOb1suqVJw+WGe3eDDszyWXOZEIyvk33tahC/Jrw5F3eXHzHqXbSndz0zMJnM78as39LnHGMSYD
dQbhxZ1h7CPzApNrJ4b2PpMijZ1/7fFA8VXbnGEYDN6cuoOZd3dS81iFD3LfHg88SiS0hmu2Yu+n
M5oUWohX5DKJBoRbQH5/JjCaAcUP7ELWtlIqyEM2TponAMzI81OuSQ5/56CCeoqdB0KtSTHe+px5
JohPgUjbqN127G5egU9Zz+EraZfjWjmiAo3jcaXIjZzptjIt2rx6faqFaHC9EUZAKy5zE+l44Y1i
lU17IhA76cLI7Bba9VLIXiPAS360ikaemAsArMa2YOHKpjOhuvCrkUhr564eamPPheuqT88r6dP0
OQKYMMcCTlftF+NJTVNRFTQfwgzENV386U9YyGHiLmJXkoYqYRaxsVp9sCgFZmsY5H9ZT5FaHt+g
AT2BBpjyFeyG7mjo0msr6RU4cMif/Lw27MGGQt9h23uPBF/mLQSnru0wnVsdy7ca6wB4DGLDPd+w
OCpFHzJELW84hYk+Et+eI033+Ux6z0WTLjS0s7Nx6TEQ+dze8cbOt2ziu9vChqZ8lglr/nZlNwNj
/R7y5yFr21MBiMoQVfPyL4Q+Y96ak1w9mGA9kCdfQ8/B00SuNvnzzlz6H5wyOh+2+/na2oEQ99s2
36M1MUZi5mGWBZhblkESXrSRs6wzsd5GwQwXM9FPbnv9Dp8RUkgOML3rY1nsBrrVC8X/1DnQqvl6
PXGye98GuqZHgA/CIubR8GiceWUnjIc3Ud3JyEqqDO6QrPeyrJSqwcMzI7ZjO5TBw0rEqE3csuhe
7rLNoB88Vs95XcpjVdiyL3E8WdWO5k/C6Yj8zNd3+o4/ihj3qkP1e+awWByJpujch80b9g7OYfWU
lcCxqI3cgeWaSdQXhovlUZYyn3Hl1/SV9SDTqWn6NmTqqgQ8Du0nxCqnAf/GWPkFqO/8H8L+gmbo
WGztypXCYR2vCDAYSkF/vMbJ0DUetTSo6Jmx/ny8rRrs/dMwsEr4m+aCik6Kal5puDGXs5WHw2x2
Lg5PVD4hxMwiL8v5wddPRaNf3H8Cux92HYFKwSHfyXHi5KCoKemHbD6ly4sMuix2n1E0t6LGoIht
etxNUC4xGpY9Q0UcTjDTKFAMJE8Gq/C4egQ9Ab5kTmLa1+oM81lT4R/HdIVJsS9j9IRVrxExddqv
LNatKk0dnGsR6Iu+RgGSIyhYtFhyKEvJksToXzK87CabT1ekNKUlYkF1QSbH6qY3mHex6DxndycH
bUmuU2sF2jcM4Tq5oQ7KsYaziOsjQ+sbSADarE6TxgeO0Y2UHk6PzQTWMASRmd88mdl7sP/WqNaQ
IJdzXmpdb7CNjwXK7YGIt1AstuhVOC+XwIymqUwllduTXz7cH/Y07fyttHfmqe3D0U78aYeFhrsZ
kz3f9lkhWfjgSxhAdnTXHF0Y62Cyh8SjWmuphxA28jatA+0Et6PNwwfs1x+ewZUirnnXzC2dIBsi
qbNfXmO3uIePIl61WIYOWwmTRX9wF4e8m/vqwO53LbJdZv2gPHxXJHEdEGAAKWxtKQJsYy5eN5gv
BWdP5yDllGmN443iBRVgoYc58Cokq5bFF3QU++8UZEvvShIV2XuXoroCdr6dFBPJPfDB31mRMbdG
pwqF58fInI0YBLL2z85z6S6OFROUU5bI/+a5l/gPla7GIIh2XvjNedsJHtIO1nxtCpbwhKTJBDKq
iVnBypmrnK/v3uhdOa5ex+4ls5HkPxfWaBXEvlXoi6qJYNjBWoFIaCpDl6vzpXZR9xeWwvm8Frgq
cpYhAVF9eW8OqFD9s37Xg0b0jjZQMx6FEI83syJxXW/xJedkPhXL8ifXzEPDNqRTsrsxiyvSIeG4
HHzH51cmk9X3Z6cB2qX010eVW72y+RpRxXK5BDEDgLT+BRquiXidlWnMdcAQrYlTMtgcgKp+dkeZ
w40qoa1IzfjImzDVK14jBm2bisxQX7NyjiIkljdIwnygG4GLfPcVEUfTxaOij3uXBImPLVu4FYz/
FXWMbSTbxg34MArz4lr/Mkics2pBnQjFdAbQfZ9+cB5DbY9C6e/YO0cFSn1aOt2K4bpWz+5mqRle
bXaAeqa33mVSkJvVrFrgfspVMadfk7uyCu9XxJMVcnCLBwS/MNxp6s44pa89Gcw5qe8Uw1mShcZe
GuMu1HiLEOOUEK/8H+HQESXLvSw3PNKuC6xovFmA4VTYl/82lCNgVv20Nphyh2ugea9g1VOC6ovL
2RWgmXTJ5yxk8OLAWWXH1q1Q4+pQ2kHtcnL/8TfzkCQZStx+HKMZ6SIlWPJ/BgwIix2H0JcAjYh2
D/gLkqDNLYXdomxKd/gCUVuNA5uHeui9cTzjZRTCbMpU6h3Od3T3Yf8yAgmGaH4ttuePRxB611/r
L7Xqw5wgzJGIdE7yuKbLTkNT/CgBXB8m4T+wOWwYeqDK/A3KGLtzORsDtpUTs/L0XNZTcpK+tWet
gS4rO7oCXZp4qfK69MBbl3iJ8ZapB0LrojyStHxgNWiNkLhPL7x9K2YEfGlEJjxxDLBEbllEdkhw
98rgrGd6njMJ9FpvGFktTbT7gvBBx51haZI74OkT9nZIUepoP0ASd7eoavvYO4J5djvKyn/hIds4
iPzYC/O0j6oLrs080P7aHyUFkS64CkhgHqxExf0sJ8zhCvimCgSsehqqORy1l3dbHVLbpdCaNvtv
JiztSD+V8JhsIInyITAiY455Uiov+YMAxM7ReLTOsBOJ5tzRPdCLZK4FJvEHBexW5YEf8FN/NJKv
f96ZllfoBRJlcT2lMGRlHYSa3jngpywsQ4ofTEKJlb4OkjkTHljk3T39/T/JC4Two0JVSDGGKVXW
YFRjaLm+9+OvXkEaYkOMpvIL2FxpaxkyU53jrOS5a3seTE6Oy31hGI0V+3KBK/DlHNBIwW9tj8Dt
IWfRiJipGrspvSe8c5+nl3UfHu8UNITG8if+lI3GHG5xdfXjRUHG0T1N8afACeHRXNlaq71CRhKz
L592RHb2g55owAzEv2BPjHx4Z9dfWruXBs9VWwPaTvuJurAqXwG0Rtz2ewn8I/JvoqRfSdWZHf9Z
18onvurgo8yU58CMC+ZXfBu4ZJzvLemXZLUXH3jbvdNQb8PQ0ffH159xlh2k/QAfhfeXOplapTR0
iyQ896y3VnIN9btVSrDUxCVNLbr0ntr262bLdYGjQioYI5arsO4dxNSglDDAHEriD2ZHuiFtMtps
b06Jw9kkj7rnjneBUCvle8iY5EyIA/+lZlByU2Ph9BMdI2Mq2bRTKlv6aLAtCm5cFH+TYtqQBJWG
7cPeUgTQIWvBKNjMQKVwhbD/aBCQsvlwzERedp3U6arHwH7751hjpxcotgQ6jkiuQMQCXEKLENtN
TqNxtLQ5hZF3J3Fp4wl4WA40N/cGeTxv/0jsJqR6C2pZLaza4FYKhFAd3dTTDIhBot4pKa3kzhXL
x1uyB31csTK0ilYD7kd68e8sjkydlfobvMUkLICLdvB1LEv0mOzm/X0p+D/iSJf6k++XeCXSIn3J
/FsptFc8enuF141lnXaVW2vrGw5MHSQbEJfqQ84aBaeXGvkuCo14QFWtrOicqYlB8dR+9lalUzTY
t7ueDmN1gJl4O3Rl4N4bkW9OftZGmPjbY8UcGy1z3BGJdHA84l5Jj3QvDYxBykxiArK23BntOgQy
DfWd0z42Bp45+/pugQjipCX6VKpflgzgXG9fgP2SsaBBBXq7wq8e4MUkIa6uOQNKDT9aGIw3HMjS
PpiSi2LK6hQcx3s7TDb+O9DCaYEOTBeUxdcnMqZkp5b26xmrDULJjHvSrF7W1Q3+vMe4W4PK0bL9
l+wMts+vdXwLRhI9a0X3Kw0MPWTjxVxVCONyrT0bRLAONhUzdUuJz2pCpOMflaEvUSdAiC//sWhW
6WOCSAMiyBy6DlpaB94YbNKzA6fz5WtyyAcPIaoxqvHaHDeB+2m+rvuULMGxNXPZN+Sv2vkc0c2t
iKeNhqZit6mRSlpen6vfbsN1rrYfnprzPl5DAUcjvcOlTnD3t2g1XZkA47dT4oEcSpwPSyLdqAvD
wKBOD1zyleRpv9j18cT7EDgnP7aviIR45HpBq+l/aVuDfl+sAhCdUGU+u41LiR3l/or7lOD2mjH+
RmRLp3Q2r3ZTXfrBfJPZbsay83lfLIDWez8UMHvwSvIZ7wzKh+RellXb+67S5M9IUdva9kuZVE8j
twrsplWiNbZgWvxvgbRa4Gn71TwD1hAYnbEDT+PGIlPrRqKkDpIoP1LB0YApd/XcBtRguJMGKci4
PGWfBVcnevzlqWFOZ+9Cy4+VCk1dj3oCPc0ARTJwSVXk7EnLpj0TsaWmGBmURD+KztYIy5Sflj2/
Hp0BawYJZN+xvQHu6a0mOVphQQ1tEoa2EfoTIlp3pTzMBJ1KnC6bdD2uG7+X+ZPeeoUOZVJdR2t3
cW+fuG5u99E8Gh10nnQo2ssv/YCJG2/cQDMswrxk1F7gAHEkTRW+Cc6flT/evdy/DtbKZy9fkdip
g6oI+buehDDPfguH4nt6wwwtIMD0+KixfnscsFhm6DFMOfX2mkxm2P5HrHB9mOwoTy1UZL86oGx+
6/vQ1DA9bq2fz5czQTgZVWNukbSegMTVIISPLxbv8YN6Mo2jntEpcY6MN6930uR85UYQawW8EkJs
HnfvbTWWrlWJ6OF7oJJVCjZmd6zHACEFG3owvkKyOR9wObQCIApOQqxL2tcxykZjVT/4Fi0b4Wv4
tWlaJ4be62iYbSnE2wEa8/wT5tACfpNEOem+Dl2ZnHuwMcKuNfMmhLiQ5zZcZXBTlfy/BbG+ezUv
/MMWTq6Cid2sGAa6fncJlH9OIuoAtyGVjbN2HzqFXq3shEuJTQkMEnfYAoxxKbMlISsrUxb0Z+1g
SOMO9bxCaa5vlScgrmxYmH5QHOxT04MpjToFej4oFm1pN9JNG+awc+AvEpj1cf6Hx+fU4UraNGfD
JFhZu9u0DoG6Wc09Jq16cNYcdkjwgqqp3B89WUb5iYMBOj42jxt2TgHPBPiSj6FISMVfKR4ANHuP
gzJn/h9XjrtxB8kaCtat3d66WxT62uJLOQzA8EDbsI6/AMdqEoDkr4t6bq6n+XWsjLqQIy4j6yLB
cl0HF/tX7L5/LXHiemFKX3hhsmzHbdekUgZZBEKSlOwWaIMg6h5Epy2H6ays9+4VXjZe3Xvo5hSX
OksoiE8bfkO+6RLfAijiLKXLRngY2aQ6ciOqRmw+ACxhFdwP81IdrNTXjY0+VEhmZFn5UaX6v1sI
JvHAaRwq6sm4/QVBlARDpFTHwiPKEctHqU/ue87BYsjHTHDXsGdnyO1+LRR0bRfopW24t+mYKV3K
Zs/Mc2/5lCwzyZrWfU6ezpD7Aq188BBn/ATaRgAnTAMJhh4I814WoVKhKhGB1oSC4GxIjaa6zEN4
yRK3Fu9U1Jei6iaU5v/SsRIZvnYUK0h6hApio5NISTF2L+jIr2as2/OEV2K+bmz35rDFqiLo5DvI
bSxWEmOreSgnolPnORIKBRleNzMMiCl5QJU+Vk+3VqkD/+vPtLTNBHGSE9cl4syiXex5eU+zi5tz
xc+fyv+n6tiewlNe990lNJ9+nQvnqLuF32V+qz1UIPx39xkdmL5WdWS9l8or4AuFiYHdT2CtWJlz
D5ciSn27kH1gSH0Z7rzkwPbV0Am+C/UgAkF4K/sSG95MEw28PUyqAPx9h9hp0g9IsZdmp5IxPqTD
XvLPOHfK8Phe1R8jb1eYOhTIDFR0RkX+wjy2WCW9JJbZ5H61Cqo+dsBQ2diwPcho3jgT2uyv3fte
gyzx77LSJoTyVF7jpu+eOFEoNcUAebgj8siG7z4Yfxes4f4bh0YlJt6yaaM/BSjFOusE3EWGz67T
vW+B+7Ji6tztfjMoUzPrRR4IAv4TZ35IgXUa/B2S/Dxp+DjFnc41thucrBMVnb531s8h6Zlk6rTl
Pp5I6q5Ne5vDH28hNzdrNjjm0oAMKmhcHIqbtdUaTMpV03Za5Y/EI/R+Yj0p/Uat4MQezkWsowYL
OLgAew/wtx/n03FB8zeFh4pPRKb89qp01RR29G+QBXA3Pd4uuUIxHhf7c+khMKKnQvgp2yTWbhnL
rPQSX/c9jzhY+DW+oH1jibDhpX6Tu0nwVGvWe8l/uYjP6hFKWMc3FLc55DzFHaZkklTiIcKJukBN
37n6byZ5iRe3sAn9tmNFwhYWSxJtQLFC5W2zwS+eC3FyywkaGjsjYlugXgJrhBo9/L+jA5MdryeI
0fUkHburhvwZBRLeDkdTf+Mvc8Z/N5K8SRKEUEEoSIijnrX5/gKzB7J11thksjm4TzeoDZh2XXQ5
gAFWjv1f7rPZInoiU8xgSWSIH3pQKJsdwumtAeWnOt3x5k8gZDi4et6LLatKJf/7qFJSBNopvh+m
F58Kd15v2NgiRKQ5045Q2W3sXUvud+8d+MZZsYkTwBpsTfybGDCOy6agBvovONcVnKpZxPn2huxn
1r+sqd6eWu2igsaxJOCeK99mLQWyS6ZPesa2NEIOnC4saC0FqPFsdq3GbKtuaSGK50xQ7VrswVGD
J3pNFop5zNKadFymuHUWm7qPqPUe7ovJWUfI1wWTEWvbpuAIaiQCC9DeOxEGd0EMswK+OxSdBPIn
I0CnC5lfL7+wzPXcaehHld9Heri+rAb228kpPMyHBi38DoLaupYpFrs5gh7wvPP6MzkqD1izolb8
pth/JD4/hT5fV+IFZUW0YJje/LApUKmCgCyaVLALxqVrjXzAfvbMQ09HbncEfZ8Mx8NfSeDSElCG
Lomms3tmqkDJH4s6kxWeE9v0lS0AWbjvIzclA+qMPH9ylKJHbW5YTGK9Bss6QuzF+t+sIXmHE58P
LmqBzuXADSSqsM3KixmIIG+S/QSmD/A6o44Vnrl7Pk/exAg+47R+P1b3XoI3mfv2dlOCjGFe0+HI
mtPQdzfdBlr4M81IjrJmn/qgcuJtsJ4pZHJVHm2f4EYAroQNqd5+EYONOt+SgLH0eycKkKVbauBb
M53lRHyeCB5HKiqhcJZ8W8UT7OUhYsNsffR1ejCVFcpyTn06G6KVgZ/+AeNHjVzzwcQIZ5gr+dEs
3bPMh2rHI+qfwzCF6CpaNQ9oh5NeE4Bf7K7dO7YMlu9hrC6ff3k8VSHVJZBWm0plw+TQOGL0mjnd
hZlyAkY4pHCg928/y/5zloVlWh8MO+A9/+MlQoZKvohTeHLEgD7LQzEFBkVX12+p4OCUeF19jh8a
wUMbQ8HmPjvzClbtHxjNpkCkPWyLYqIVFKYcMuCNSi5NfeQQhSK5eaKDxkZurP0M8DtVpwPYYjgH
uMdQnjY/5zXObjNm6GriWI3TbiDWN97PrzmaOz/3zTh2czhjV4zsKPcz6paqAXfab76C5mPZlC6Y
eEjJMSM3+0OaMzTwttvXO/fCescGoQPpXvglM9XePhM3KTVilskP1Zaa8TlSKWfrn+ushYXNk396
IV/H4WQ715+1pSo1qQCSQ55+sFNMpSlWwMCTiRb1tP+pInPVFnfJnXl8ojL/s4xLa0cUwKGyST/6
Ea56HJofxW4U2QTW0g1iZWx69CKKPmcm65g9/aPAr7DtNx1CBs0AiIXoakjVCBBZpmgX9AzyPS4o
zxAZV79Iju3R20kaIk2gVrnRslm//NfX+aHe4e5QGY8qT3gpJ6mVjoz/c6aTSWUBy1ApAGAEFH5t
Hr53icik051/IHBFZ98sSX/1fWZTthQht2NGkz96F351/D2xoxNh/98x0WCFDl2ia0Fdd3cvLiDJ
ZvX/NbCRLFmMfCFCENChWLZzyLsrzrlVqOrhW9KOh5nVovMddNcsbasjiVVDy9kBv4fP5uBxUZUf
N1zrOSJIJwRKMy4kj1QbFykQ54lomkLZg2bcsJnnuvneU+m2cJFgOfKDHsh15dIRtikthvN+PHSl
CH82uC/D8tJWSWI91VsfHORrMOQyMu03IZioH/0jVeGd5mCHrEWL3IOX5dXoQNwmRyvOhltMNT7Z
miuZxeiZDTjNIaw7Ab140l0VEIt6ZKJfIOesX3V0MyjyZZR4egSweLvQrgstHiPeqy3FYdzC6ZGj
nMa6y1WKBVVVI7UFlJaHU75x0QEWtNarg57MO6HIFMk1ZYgvdguenTrBunvHy7yML25RNwaMuprp
6H7T5BE2NenWKg2ewMI8/RBL7cR+7VVzCTgtyJRz4oVcEv3+iYfbQ3IFCDpGn3nC/gtjspVsVDNu
dP9StSTiQgr9QoFkHjITaHf14Bx+g8L2rfBV/aXUIbngCYVEy6FuWp8DthKYltlOk7/FRnqYSGjT
kw3b9/BwS6cyg0wyttmeCZ4DNMVx56024sbgVdJ/TjG7scpQzZrhHVmiIiOnOyVLMOasts9+WkEM
WyXKXUAfy5H1Pmd7K0FvvmYWvdTFweAiLRNQUMovgWOIY4fO//qF/ASERX/M+g9UbyTBvz2ERDQu
geGYdAriSMiw4qQlupcmQHW+lk5lV3q1i+mf2yPtAOP28gzpcpYuA7YRh0zYYA7ID4GDbOkVM0yT
fy5INUqWC8jXx02Tb1KRJV13O/mwsiujny5mYNlIf/HJwyj785vi3T1x3QHxXCY1764xJOLCnIJY
TRFs+PxJwoBJhMOKirK9q1un71D29j1+UhjGkZUXFvnvQGu2+y/kaGvfGvGhOTnFhPBiFtC0dY1I
DL9ZoACheBlwCLCOMFdErcGuNkNUiZYGLhfSZn3pW2dEiihYmQpTJvTed+oflESDxIwClhVj+KNl
kN2E+DIC4/j73JZVwd5SrSd0woWx13kFPzAzr8RDJCJNoegAXL5IKitZ+YZJ8zMTE8rtvBsGN9BP
ttyuuxaSNLR+e1LM6kMWUsaiJQ5guGA+wCqCq2jEHGDUBG9WKebJwX30Yfn9CZsaO42jOTRmH0DE
buZS+vMTuvTvfmJU7w2NDPfvYDBCGLTK/E3NgtukJ8OVCjeiVHjIDQzcfvCUILf3dugw7MfusIME
XRjXa7Jx3TKS5FSOstuC9fHTj7zmvwDFF/xRxwc9yGtQLH5kr0XpIcPv8Lxjs+m827SLubE9jW43
qaMv3LYhMwzuLBLClA7GUx0MT/+IJmg6+ZNPOO/QANh/JS8fdY+9FAjLGNZAzrIRtmHUJLOfJ/Uu
JMsPQ1F3I4tsafiYL2hFgUGe43LtHF7fXB26TNYWDFZnrDAgGdF8Xvxsr2hjImUzPzKAEvBq+JiW
jl+N3cnRnbm/vvadtONlLfmc4A2vCUoauf+FckDSlaXeJU/p0ChmaFjjuhVctCaPWfXaJs2w/qFY
MLjRlT8aNf8jEKry+fLLnNK2BRG06AuQt6owGWQenm2ouNWFXofBeFaX9tXN3z/07AKtH1m2JH5/
5eTOyQQcl+Hpc9R0d9uBF39WeKWsZunejoCNDNPZBsGOu+TEZT4aNcTM6/3+5vRj3tFBZ+H955bb
Q03jd4cmlSH0agRFxEfAykpDqJbN+j4JqpkAF6aY+OOqO/e2nO1fuArBuUzzaxYEuwLxJW3xoR55
TuNDLHolJHDVhT/menz17PTRPlGSNu8N3Obw37pQL7xnrwJqOWmBMwfzMpD1m+saQtfd3VSfkw7k
3cPLiwIAh9eGnDX1B82JcEbfgUoKmunBFldTWqvsIrjQDWtvBAQuMMpdZeKZ2FstUU4AHHyyJWp7
jmzlqXJTuCvhUopQRtsBnNbC37qBm5LOdWWnYIHZD/nPaLsv5upV/Lw1o9FxEz7iwZhSzCEwOGgi
2hIs6PGwRzEaXrJVsZ3wF8PaRivhTvACJic3wbD5NlWf8fq65R1O4okC9QAx5sUHB8vbLMzqcTwY
M4jXA0LU6Eyi/oOANWO+3qj0e9PvMZDgKs64Yz+K/TEuz78Z/tVSz7aiTNpBb4nGWJgtlOGZbsHF
D76xhSDcQjl4XJ4V5Yn+5oEWKMAX6lzLRXOUFug/jv9gkcEH0i7UDqNc3plXDilEBiA5T40f5yG+
N+4y8tMbcjLhIN1C99vhHew7uFrQli48a7e04293uQAPkc1GH9IAYthAya8uInMp/y7TqoFc3YoO
MAIy1hrYR0wuMLo/R0gDIH5zxL4QHnACh52YP41i+vEMCsG37i4eY/akmjaJ90OSCs3i4a8wHh/Z
UWL6+2e1Llfq7AKQTiJyI+u2n33bcSNEpFtGYXcfd30M4zW6N/F+5Nw8tpRYd9C4aI1DElYiZlf7
1oMd4gP3eBkDiwxyohtqkrDc96MVvB4HfV/HAjI1je+oZYisY5JQRpVJMerPgUyBWq2RkvofIg6Z
4ni04L6pBPiEwWCwPGAtj5FHgDV0tFBrBjFFMWkcUoGjdZI3IAIv9HHR73UsJDKytiBYF1eDq3TG
wXC7+Nt3jBsQVAqU893KjHayJTmSCx7eFWPlczArYCD3b9HqEQ2O+TPvHFJkbvhQi/tg1YoiK2YH
F0pLdtsxR8Z0rGntrtbgEsKYKbpoDSWXUWUnQv0laklekMlHUIAgmhmNOMyzPTt6c9tzg3HGbxTL
e1PR9fWgoWezgbfidv1o2s5URKkQ3dQNe0HpJ7ctkdL5h8i74D3saHkYc1NaLEomRjRgH4DUZAzp
WJwPHIjOLtVxMBxSJh84KttR/4S6vDviMSRPSccQB8+cGS+gD6GU9MTR6Nc16twrD2yBE3Erosy6
OM7f+SwX3ADovykNXPma+EcapXDYR/7tSmLc631DU+8i8LG4GZo2pQJFBAwaE/M9Wq8g30hhqOri
5kSa78OwZt9i+IebiaxaEm6xU4Md23d8lJlYpn850NChXFJj4ygbhFKsMpNo0m68XxQ+XbZm3ed7
Cyt17SQElqMVkzwLVN+0OcyY7GhPvbTyI3iOyuBlVYtKroVMEz6Se9QccI/0EBBwM7nZfiBQAGq/
dRHztqCbPoj4JXPEKzfOU8pb6YDC2bJen+6zjZim8u22kpHYhfbKFFLNSEUmAzMM7078wC1lXkkt
XFmncJLZsibqisPyKIIsdUJQeNOZpKQh5P3qzZ6G+TiXPOOk3zw3n6zYPST9lvWcg+NQzPMDjh7E
kUagI5fkDfqgkQCZxcqZCy1GTyXhWYBF14ukawyMfew/L0nk/6lik5VJsHY0ymKrfRelk9qJ4qHG
o1sZTbvMl+rm5eYiRIgvxKOcxvwZrDDxKpfs2qkjHrwOYM5jfituPfsHr3TJ8SzpMmdC7Bsve6bc
+GBB84ad+9LWHVZiDcVTpAofQ8MF0vSdIxrgGj+8TaXrS6QbQ+JMhJORSWF6bHdJd2Ki6ijU4g3G
K4M1WYuuMABRrj62vvzOAlv4Id2o/ykSQqCcQBw16Xy4H8wHC2WUl5S2led388/BoDzSVxXBIOu8
Z2shtieZWftBHoH0lBKq/5j5fe+MzLHiqemMuekDzEgXdX2yrD0XD2DZZew7UoWOVlZWUTmx/5Of
jkJvQJ+e/o/C+tZhSYCOfNyapTsFHGMj6vEKnSlBN5g58ruBT96vE73CqIeKuo4rxEWYhSuq+Ct4
OaNz0TyF+FumGGK/0VImEiyCP1su5aCwWG+1igkEBwAoV9lkeOZrudHGw1fquTygHk9EyyVW7IHy
i2a+tqe5QPEwZ2U1Fn3uCCRFBdOzeItHsNlVxPMPr5PSGE//0EDnH9Cb2dyLVulLfp3RfyQeF2DW
pk93E1wCKCYlULFeA3jIkQOORihwZvcrE/Y3xNQMf/LFbDLgvcFgDVlCndDwRa4Kzntzx1wkJc8R
1m+GjnCNUfcw4ecWDeOSiz4KJC4y3FEXP/+5j7Frd7W4VbWAHvmzwIzhkvXT1Pngih7JPB52zX70
DFERUa9xPFi4oVjCiDEphqkfRftCjpnSLIwRD2oFTmPEoYq2NSHhHuEpj4UlKhmCsYHrF4xtRhHn
POVBhctVMlp5IOR8kycUWFb6ATwY2BqLhzKWNHSNi6wG9JLUrfRXDvyMHrCGAuMvt1dQijusDJ0M
nzJ4jZ1rM0WDo/063PAs7cDTZtleER7M5elEW0gUNAoF6Zb8fOxwqOb8DpCXJLzTtRbiKuDT4Sfl
ir2PuOLLK/8t4+1JzxPzJzYVfUoT0ePYLD2IHCFRisUYQKzsW6Ml2l0OkkCrLjCghimHzYQQcsEY
1kDbmIJp77uvEdKo7jSbVq8XAckcWvqCrLiUEC8ed9MFgisHa5zoJBO/PO4zzAW5WYmjQRerxlD4
gktWH00Ca0nnyEZhaHyQIV8sH6x+1dl3JUVm2GdlvcNVc46b2YQjCsjL868iDu6+VSM0fPJUzhB3
7LCXudJpY5y6rHO2hGnoO+1gDsHCVUgCq3UDqxqPfons5X+yuaLZmtsVKfQgUItpGSSVg9ZV1zrW
FsEbFilzg9wpawQ+qwxicldIPPGofbpCZAA5OxasFAEU+KqkQzW5MhXobz+5yBSDkxNZ8owmU1N+
0R+tKcNQBSLQjdhkRjs38ssfHzNZRPEM2ZVPCALJISP1miYp5AVi/36+UWN6VWosxtFrOIKFbn3M
kgabQwVwQNgESbbI1YW4QJ/YDkuJLfYgXUus5ajSv/uc8a0frrTW0lW5NZLiJM5Mpth9rVFg/M1L
z9/S5wMOGWE1yZLh2m0PV4C6jr+0FV8ABH2jFckd+R/BQnybTZ5LorVNqTjKS9sv/SLY3NpIYrq7
JQF3J/fLv+9lI6D0XIgn2231cFGKb+F7gOn34cKPW6wKvAs+g3ffUPt4eCr68MFynR1XnJG6Fpm/
q/k2pzfJDAMuKITpZv/RrWlwCTaCeNVA7p3LnXe39mKzP0LNAqa9Rl3tsaGwubW9R6PX78eIQelS
jzkmtjLd7AfDOXkf7Yf8uLa+GAnT9FJKmQA1ja2AOfN4hLMvPcme6D53vPbA3vm9JLSx/xJRoYmI
IzRlIMlX9U9ZeX1uAkLstqqr8BzcSLbtWTcWyNd9wds6NykNk8cxvB53jIPIJIQnPzNF+GI1tXi2
SjM4fNKg3t71oZzHlTdd1rwv9HIZE6mtT8kQNZu18kNNx1ne2o5xSAK2OaovFYc7hs9w5UxPZlYx
Mq9YZw1GnsWtF2+eCNz2M+ArZ47f9HdDg2AZK2nFcXjriPme2RnB9c6Fi0Kvv6wNBLA1+EQNDWC8
023f6oFcTfaISkHS27hIDcPVhEkeKeU1VvRrvbgPT46GIL5KANQjU3SnLKdpYea23f8tpoJdBojU
Q/pYlSacIVHE16xgxRBEdV/dcVveK+sZVGLgU7+hLoRybva4YlFXcAQ4JYrkTaJeNbTmT6qyUIC5
RleVUSpR3Ah7a20fBkawbGW9dxzmBs14hwut86gHuDhtiQYLxnORVH13RBwumbdTF7dCfQLqnpm5
Rq0gZpUqJocEcwi4lsOFVvfQRUBC74zAxQAl/IW5CVKSGXjUKmF4h6kSTgK5RGqG7P2SI0D+W8B/
4L9p27/RCFqiY3Dvqs49RZgne4dFNne3dgKgwwA8g4eESYpdgLuiElB5EmQy90LyguC5O9GInT0V
P8Hddw2MCeSbxgJon1XMMO4YX9Mb130Pou+mFqb+yEyPds5bMBHxlQkHDugOGnOxwLH1iEqSQ7ri
y6Tsd2EGAZ7YfBtz5Yk7ZecE8zc0j/T5fLZV1jPbfoxnLDKyqvCezNwZ9tu6CHoc89slys/u+Ac1
JJ1lQyqz2T4D8jp/2dZpPboMka933Af33b30e2YXbUQS+5hdrA7j8k5jtpSIHLPHiHHYxzmkuQ42
4JCPge1/iWx5r1mVLXT7fZS5PlnKZ0dVb9QT3EFNSEYX5AOxyAwx1Udgrdc/aVShJZcc4ck94OsR
R9aBJn1MLCNZSeizfHUEyN5NYdrxAbx/At9H98lrOaJPErmqxAPkL/vij5Sm8ZzgPXgLIyXq1rFi
+phHye3qOvOLr7QZWX847k9cix2AWkgaG3Mvhwp4A+LeIknrs6l2fz2lj73sNDr8RVxUnAER2XEd
EWLIUURdMTY245J3acDl6HS/0tYy9COaA/HsacDlvkRa0vAuggbNYiEZQhLcIYSMnWeU3N3FQ8EF
tkii5V0Se2RTzFJKG7XbZbaMw79m5o1DSfCF/xGtsmfBfM/jTTUzvjaO+bwzTGeAq3v/56zMFxJa
Fm0eRsxWk8cuNqH4PB1xpQhlbiADGDolZO+bZfNw5nC51P48uoHXnwXMS9U+7Osmz7XtIwDE6zUm
sH+bxemfajRPlGXYtWtoRsS0bpDoGwrhiFFGBs3JpdlQML/vSqqtg5qgjHmqlORiAdRH3gkmrlFM
RD9z9qtWGn524D6EQeygnxPyNPvVt541GFOdRew3Fl+J5YqhMKzPrLZheLl2CIfQrA99d2oVy2ky
Gox4blinuhspsMUq1ucGhXM+YS05fGDJxcq+0yBihyzxTK48Pq+qseSrT58yNThSOp9X6bg/8YCW
B5jkw1MFl0n7FVzbv2SSHxsPL4v7D7nHuoxuDgWAnAIVtKzGp7M7jl/Y+W9i43aWxHAVIRXF9Tvs
4aOswxtD/t7pVRgxA0zcA32WcZL79mRTa/51a5KkQM8xZoxpljKAWGLcPrVLVNyOBR4/S1QBfydS
EB/XISlwwzGcvtXCX7uoMYnu7RHjPgfsT0M+phs3SZTD+T1fAPVQm2U8IBH+PrPjqn+oYyfN7UjJ
cOrJ4LoWxPzIX91Xv7lnxhaeLwGNKCH3TBvL6x9ajTj31d/JH7+V7BlYdoKQGI7QeyXD/leWEjs/
AGInzcmZhB5kKyAZzb3GIbUhMblo3OR9/h+jPJMrVkVJsmQ45Eb78xs6qr0q3v8rfHjj84/RG9y+
MyYZX5G6y69aBSWx8JJIp+u1u6WiMUJ37MoJm8L32YhRKeeoqYJSwu5WRpiYQZQZjEY4Sh3AqCaa
V7dCehudwP8yEBJyB5tmHPA59bm7NEJfnG00kadfn8fKis/cVQZ8Ef4NKtbpueJ/dJR/U6Q56nh5
McRcKp5engXIF3V6RgJ0SAo29lBkfJroCzp+FgUqYOJ748/x5YUtB9GdhbwndDNJnmd/su0YRQGt
duGhY1GFsOGH1wvG2LTWDdzEc5biQvUZZ4VHgBIJC4r12j7Hm+Uf43la+jnX5VprnZDYL2c8XHTP
pHq2e7kLg9C57cm+A0mTt1ZMvXFtulNMVaBsU/qeOFuPuiZ38pNZFbx7EgNs7TRtXXUCRIVW+FYL
ssI3azhShLM2Jj9whveSMd/OmI7B2SsYqLbHbPULRGrDUL4eW6Am0+LIyWJuj1XYxUxdxxyX7QMl
FdK2OblHaTT7PbCI8B0wzeSLKysu05l/5n9ASfy1vU5v0YLStR87XIpyIWCKi5UOXsaTdW1eS98t
dJmerxTz0yv4ghl1y0LHNM1Lc1wi2hc1qUAF7+L0KQLELXHbLG+0m9O6eJtNjG/rJFLAzrGExYDI
WTJHKuOjDWJIESLnOSp2bS+9AsC8pGj+Xr0VNTnBGKzfO6i82z8u1QlUV0vdIxy7CywN1p+5SYxU
Ndyheddy7X97oSw2RUwpu0OzGlrPBIOS5uaH8Tl+7+HzGOtFBww/OCXpLkP09i+4LzYXqKDrvWnk
NjSTNpNU/UwOvIwGi7Cn4NPae50f4Vt31s1SI0LsR3fuHyBwiUqgjzQjP2kCmn+V0qYsuYJcYhmH
GXSPsa4+Gt4TMFzPfgu/Vp88M4FbGx3hfahqv44TXbdLFrSvUVWWNN/1yKF4QeKxwHt7EDIUSyG+
9f4xjJzxKNf45E3OK/vvp4SA1tiqBAt0Q6R3bwlpG4XNRK000zBK1j6/lh9DHSacxpW1r9mCY17w
cEwJS+3B78MZR3jyWDcr5rrg7wqqzNispp8Ti4YKWRq1P3Jej4F0tTLD+vU0nIFxI9EC14DSKclg
l80lZhyg5lVT1q48+x3FThPtP2Bn8TsKddCJg9wt96RE8e85usI8bVpL8vNleHoYOHcJ+O383wtP
ox7u3sxFeFThPuxTO2238GLCnrQdQUAD+9/QehJZXU9YfdrR+AR8LDBiGaHugsdYXPs5o0D7sGTA
pYri7GOoPkq4ZsttsMKwNjuvxHRBDV0yxhWIIxfA7CGEd1OMfcgWirfJu6dofHrLwx8fMqoQErPi
RNFOP3HFV4o+ez7FNo7RBm2VIzl3rJ4gnMdDjSJptOopcAM+ciET4cdBU5oUIyM/nTops7K8ixr2
AET0AJWviOxd8Gb0NZ7CNZFI+fLN3K+dmsGVQfUvUl+ShodfN8re52BZ4Uxc8eAynpov9in1u0ES
JA+Ar9kPE8tDGY1fR4Y/cGKT6pbdtURSRtMBe9H2+G8GY4jAS2RGYzW1XwNoN0xi3d6oOCUE3e+w
52fHkGkEE3xepdgZmaFL91lVJskt4fCFco67PvjGZoERNrmsH0SrUPYO36ixrdGwdQxcUizY2Hih
FvgNsx4ljIwyha1QucMB48xo16N6B0+2ENzI6moPYBpMfmAqvXeTezJWt5T8xAnJWpGI7aqMEjWG
sJ+zgUqZXofeVwGKfwhy0ewx7QXC+v4791top4CMYf5EPlz59afZQdC4Cy0dtL66YPorguZZ93ZG
+nrIYD3bOytocFE+k8N9Vf091cecwPngO/4ykvoFq7NRwnLLcqpdgcbuu3t2Tp9rTU2iY8kUW7m7
IOhjWv+Hgx78A6/lMAtGNAWXIvy//2VUO2+Y2/6whHIpgmlStv6L/Zy/Z/ZB/p66/HhGS7p/ohYQ
0fHABytCW9rDYdK2mlSRNc275a/DeiCCcuJHol9ebnehCcuJo9yXSa25k9ESXmQwdPaH77s7yCqV
nAYbkPOab/iGcBwVxu78BtDL0G+wUTQ52b2QEPln7JvHdsj87tG2YLv4UAxdRdMRXHYzwJ81tHXc
86shSIf/kLyQz1b+Ss0X/B5Y7t1eWiQYflVKQlRrUuSz7x94yEgIvv1Q7+wrEGPRYyjkdmiNPcGf
5LUp9C3Z6aU3Ms+dgy2EwUOCa+uNzQgz4g3CaKooyCDeRr/F++YxqfXkROiD/bakqEKdnFnx0QXZ
HBLX+0C3c3xAet0hrNeJl4VeAn+/eS1vos/ChrLLxxIFPj5YrNdYGLpE7blokdbGeqRMhcJXQ1/Z
hAvyaOBF0Yqkx2x3GlLeuNvy0r8VOQ6T9Xueg/N6LSBuWccsdWTWTKK7kLA79g32WeD52prBYlo1
pXKFjNB0PO1O8RUJ5HeVig1uITEc1PIT6hwGsyDrEAazoKwSOOGeLM/JBhnHf2CozoePAArha0IM
vv/ji9YgYBmAZJpVvHl7zuu/usVmJvP1Upobzk2VO1VE2J/i7IbT6dGyiTih4omKDJnVjvtot8cp
0t/m0mUnV/oA3wkqpKs6ENOuFqQPLi0bqGG6PLgGG7Gs4ozEi38PWOnr3KAr8Ff33qXMYHrHP24F
Bv7DVQwKu7bIvjdVd0S4xJEkUqdsn/MIMSckzD+7b6zICl8HsfVvakxWQ4a7+V2ZWS1j+4+WebVX
35R1USZ9rREWO2trHSNu2E13TkDBb/suKMEbBWQMVJzhaE0PFrK0/qeexlu9uAW2pq7UF2Ahg4PP
h6fcapnDuormrsUmSaU59f2TonZ7XTtRkdEc1FRuBn+TUuFDDQ6mFIGmRhjIkg7etDHvZgj7wljo
kUfWA81JRItAL35+X0HOKiSoHsgeQ5I3hjWqNCXioQEGOIpdB1vBpj4U4iMwdusIk5Qsr6cBG/GA
tTG1Jyx0Pg11o5PB5oqikbscK9vajGvK6To5zqUtQiKvWN+EJ8aieyiG4Frk4Un45SW502Z3S/lt
pymS/Gi5koWexL6+/E4z7QenhOP8b4hRWCzmoLG6YMNix427qKjD3EHRYpdhlYdisQKzTkZyGAE+
vuGAD2QRqtpGlIGvUwRzGgSgJUpTra0XDZNNVaHSm3x+jWd1LiKkgvVpt2n5Tw4y4v/B7vArkCts
iZ1CJymUrw7L6m0TLMKydDW3dfa2i6fojE/By785LNEsZ0TWEcjabTwaxfStP5/Wk1KkPDFbtE9p
zu48jmyvlMJEw2AEIGLGtik1dWRt5yYhwNqKiCCBI41PNMbVxw/kYzTDAmnNC+vuBq7V7kA1D9yv
uA1lIFKwOb29oi0fW/5NsDbluRWFIpF2DokRytqOoIvCFEBwQf7W6+B72DZfJg+2cD8wcsyr3RWw
9Jr61Sc/GvV+1Vzgg8u+if2g8sN3Bcay5eZE9zdfAb6eAB8Yf59LHms/n9CMgKlvXlxJh5dABpqr
b575+SvJlq3e6dzo3aJV5GkYMDTGLDEetqeN2xOixnO15k3RuSrZ4i8C/lhZkisIGpA1LCwclHgL
fzpNGBHEsUNVi7rir94KcnECaKFcaVXbWkGmDuFxKtMiWsNebkO5jqRYEbsJLRG0sp8Vr/5v+xPG
oBg7b+8+jPsT37aXYwg5Na+aCBu0IBtm1+04Yy7tR1yBtUi4gmeuS1dfNpCai/zJTp5Jd8S65Veb
odGykwqVWTH7cx2+8VI4r5Eemak3tCPPboI2bgcxTGr7040V4nJ3bBMDGaaGFfEtK3DEjqlI2J1v
R+r5Fi5g3xuI0MtcDHH60Mvtr8aPoQlSnZViP6bCTJSJgIbVb2tmbAZJymVb4og79xlhF7626qzX
P/J4ivJT4LIUyWRRkwGEENZE1Z3ECanMyX64H2ROGq0mx761YVIbY7IuqRIJPdIl0sXqUBz+67dE
0qIVnhxUvhJNAgzLgCBpvrfyhjStjugs0SG4IQdPEPQuPncXDNMKas40vcvm67b/rteklXeSxBp6
mozTVAJQz6IEFZUM1aTdAWTrL7wCLtRfqkfuoK6Zc/9facf/GdlSQZ7LXYapXVvWzlXAjPDdfTQ/
4eBfqUi7k/oZa+hUjVIS6jJGpuBSVgS1mwAL62naQyC56pfQL9LFrOAh7ijkuFcRPKrbwaXj99VQ
dzt3v7YlPfib3SXQTFiCjlpumIhxhvDGU4rjoWTo/zlBAsqHDhwUWWJMhRVU8zqP4Mp4h+DJ9Qmo
vcaC74LIYm6t5/klLielmlVgrkXKX7INxHBQzqIjAkgnuWx3ugpW12Xx9dfRjKvFgg+Y4xNX3KaH
8HntNAEeAOxxGq0Bstb05BIj2t2QfZmQXTsl2g1jSng+lHlJP9vsODUK0WvQmsBY0Bdsniq3J+fB
TdOcurY6u7ST4Ty1qbem0qW3wihtyIRs2CeIIjyRmS//sP8mNCVCzkLbxpl4venygExZP4lxJGtf
rbOkwkxwtLw5Bpn8V5JeWyw+OryeqXVHFY7ZJ3jKOViwBZ1WaPpKDOpLT+tBDehS1nfMbmatq5tV
Mkqap/Hg6LRt1TPA0G8rAH/Fx7wSgLOk6JXlkK7DpNRQzJzZm+AZSn9jp6XfXBakf3vpb/kMkPU0
nc7zUf8VdfMVinPmi8Mf+3Zg9Beej6nTKMpBRyRns1Xe0il49ln1ifVs7J4xq4sN0zaU1Wx/Zd5r
E6aqfcvDQQqLLDe2A4F2CVQGNrAB3vUghqKVlBN2qR5GNGbWM7YeIBzZ0LTfJ/rkEnjSg3hTxS8J
a3APk5QVrUHiTL7mObBJtjy6g7odt//BsoVRESpW2IKXqtj9udA1B2pXZhLXwbGBYeDK5QwXe+m6
hw8V391oBbdwfWohJ5fKRh4Gg9+baFndwpGULrZBgOx10m1eq2MxlQTvYeeLumFPnR2vDq72Myic
+pcc0S50U/km+bv8LjnmE3k1OpG2pwDtvnhbwg75nJN6MMXZzTAeqbOWGU/id6ZXSAuxXEPIADOi
YReXgO9jwT7ris8D1Fp/hmJG2J8Z9OAohEJjRyHr6HaVDQXOPMxA3NArHS2HkmJmR+/llEDPk0AW
XTfODGmBBG59ZqYQT7dw13UoxBxOgSbaV9C+ceE8UXE8fOJw6BdTGM9+ulh0H68L4WIGUkglfIo0
lBpcp+eM3ERiiPvo6y/qXmG2w3rcBjcl+KSUJYlzVYHvpA56hCimCCWpxRfJrEjtDN9HnHv30515
xPwTX5DzJQwH9EdzsFlQuuHT7Rl1qyiqjv7VA5T/RUuTDj2MrftecborWzJMW8F4/eRq/a60o2A/
Ble9xYd3LdDQ/wW7eUweCxvXGFfWhzHtSsqXbNEuwtPrtOi8YkoFm2u/Nl5mQxS2yhKun5bEAhMw
iWTUIaw4UeYTjFggpV/UeJDL2jOlnCyRjfYtikDQo6XkXOg/5WKGA/FXNcuaMbsMhaHO5XX3fluw
3TOQ+c+04ilSnXl2dRdKkrIxMeX6bHPy7JmTP5+ypHGVmhRWTc2RheQrO2rJmD1KF25c18DVliGG
+LRP8+WOPKH+pYJNkxrIZy8dJfP611yGxRfhGNEbZn1Au4U1xLlnVbXvbaBGL1jZFvN45GzDlfXw
Nfn/SoY2B/p4kRmMxuktvx2I7hU6BkEZxQ/GqwDqQhYUAYrniPGZ2WBhsb2Los26RTPrb4Ek7f6D
8+pJgEFCSuSqCeBea0MVqC+TfXfsQFjZfRflcNrcnuVPvkkB8AJ8WX/87DR+UZwS2zzeM7mY08OS
Otu4YTuv0rgELhH//ccgIDucvgW6Ujttr43xMepE6oKUZcqy0WHFn6SkcjQ6wORuFNDjggGLsgt0
KUCmI611U2QWGTUm2UREpaDgnyMvDetXONAKNjowXGlqUJykpwizI1FhKmZD4ut20sRS5TluY/Vi
jgr/RrDHZD5CNvGsa9V68SUWwc1ltLpTGM9Gq15UEYuqlYkGr2gHL3PxzxtUkFcMZIvculfJLtQS
rpKpe7KzFJ9WM6Z5ihlo1rQI5SPRTQFbLKfptxa+7MgsRj0vuxJgUhtZDNQ0vqufP0p5Kj8iFwTb
1ZGRHcwxonw0qQmO6iJG7yXuakNYroiqlIUVkPXNgKamyX/B/ljwrvY6O+XCP7F+uy+V8CPOm+lI
J++tZG0nMmpcTkdaWREICWdJl9JDHPqzRtEam0F9Zrj4nVRFITZBe0jHzG586xSnFLcVBZoLVpve
JvYZnVFX9PGrCTEbIwFliavCVqROLbOg1OxkfyIXrCpFrSAhQMqKvq8Xp1stCDjzECWUjuaVruSb
EPayaD/pXNzqdLoMsHys2yKyb68ywWtxUeMlN/qWqGgoZP7fzD5DRVIV74+cy5Cg46Mn4XLy2HQ9
zeTtij+AuH7ixfEkANmls3+XHpPidDdR2147DcuBOKdixePGmrIfikjLasr0G38uMudA5vQVTzLm
kMJSOV2S9ejBFJZr1cQi11yDGxtotEuwtXrbeCTCP2LGy+SV25vap5cPzEatzDgCItZGeWxLQ/r2
RYJkfWFevIzsQC+/xro3tjhym8cxRf7FqU66mh9kHQTa3PFk2cipPzlaHvClapHdGlQ+7rdO2o8u
4JRB+QAHOw+Tv5z0HaIzELNKKk0+KrCBIB4LegPtaHP8GwObnkW6AmbrE+xgUc/Rls6Ye9XbdopB
8LYaCg+ZS/uLXGrhXPrnhKU+h65i8Omf7kk5JAqjK4zglQEi1ONr6rTwFRzDGwZNpPpXCEVOcLPh
S+S1KIe4Om6L+rwQTx2rNnsl5jOIInDZ3dKwyGC9XiMTBsJAoDChSwRFgqc8CATScE9x5Edl74yN
QZFy53azrwpmPrS92WrekkpHqlZtN77cZfFZ/BkoiRDpZUx78f0N7d/KIUqLqTysvxFf+zlrcSMc
uykH/empiGuRToc5k2lQnnaW0p0pBY/vHBf8WkriuA7URyzq4zuhzWrNrEmaStovUEYWC/qcraeu
h2sUrtGAnhOvaBY/LbFy1w9ZgCDJZAQoD4LoiByMT/Q4kIx4cPiMlnG5He200WpUpu4xsrT7wB5j
usAdUAoczCMcfVA3kFZhdLbOQJfCwOZVzPOfDudwNX6EynHqY8KDwi9BOKyr/GooCi2lfPyqcRdg
9pNskkYKfO6ej5AKBSVVYw3rjo+XqE2D43fyZk7El3wkjJ1CvQq77ksrSliw4XU0J4CBwi0U4k/q
tfopg8Q+MyjHPj7UX/WKMja5b8P4iFj6LAOqR+WzTT+4/zuiAq55/5Zybq/F/LI2JTPrCAtJ0UAs
w/pM841V+VY6ubnzjA/xCvBU4bTiGNTW1/IweACrQEevYN523E0sSCVtsMlKbFKRVI24N2+WDJsG
u4kPNnI3cgxvnsfVKNERxeKFExdSSeNfoDbYKvoAhrPXIN6xcE5RA1HymBlRh9dXl1EPqpQZJ/qZ
AzJMSDuQEC7fpN7haX4YMNYAO4SG/6pRf77lXZ/DfLBKh4kkQxkqlg0LV19BHF0DkEOpqYJLRC5L
oWObzN7s0vwt/g8Sgtu1N6YlMNp7xXIjcDknUHD6yc7h2Y1vrudwPwK1wAC/mDYi4UG5UPLCBBBm
cbXbIkbGM4SWb/2REAe4W11gGVfnIYFvSJ9WY8q2u0nVeB/j4r/WG+oDBNbgctTDGgP7Bspuk0T3
/tJNPuZXtPg4fHvCHtO5M8MhUuCAF+0yOltivuHVVS3KGn/BgWNRUQ/gdk1sbJlCJiTqu8zE5EXf
SCckSqunYSXzEcbyrs7QmP9HWfZTLfDYDHkLemipnrfQB3GoQir7Y/13HSBV5AWukXW0/m8px4XD
Vp2dY/MXbrOlZY1PvyJLUD0ds+aU9GRhAs/DAP3J2tSdlBlU/kOoSZOyg1wgaXxNrrW982gByrLG
yXCS5D2Rp1mxc6CA//gyWPrIErR2hb7uC80wjNOwVReOSHZHholyt1PcoNDL6RyOGJUN9J6Sb0MO
nLLLqdq1BTY3Ol3eyVJ5d1pYlBP3JZHNuJuj5zofp2hhEq6PoQ8O/xHPSIsQWUp3xrddS/5QPm8h
4cCyB8dIZAv8/jVonxAwn2KUS0eMksgOtOANTiBMfh5iEgl1YdhzmyzWuHeQoQFmxD1BGeS3tqJh
7M8bDeQCfZDKz6/yU/t2F28NpE/g5FiuAkiyTpBaFaRWdn4ceDtEoVXYfwr2ybKLnUsEU/hbGbsQ
LoRN2DvITIdnuoLBqzQgXhpaEsyN2h4RDxzr+IENG26ZuTg0w4EaV5Qso5hAPUmEX3/P2EgfnKGL
ucky4m0T9+vIWKLGpNzzaeoiyBVxEZuWhqKE9U+TiCHcKNIwU+UkThKaz2sTUJCrS0YJ+qUWtIm8
MlDkvz0Xcyk1QeGM0N2TUYxit89G1pk4tbeC5V+IR/fAGavqejnvR6P6L/mD4pD/sBxZwowNLc7D
EXy2XipLQN1BY+uV9F+N+c1z0U/bp0FUcG/Ln7SU3XFPvbuakbXVeVOii5CyZWQ+bCZI6HzyQkQk
j8JvulX9aK1XbcR4fUuo8ogjvccZdDbjbwwzUPLrtYDCjOxfrcQaVlQ3LJatX3SsPNLQG9XSqwsS
9dVAsn4kVBbFEy4eM/twGL9zhlGO46Qd+XzOBjB867oiFJ3PqMa1oPtIsEBNT6Y0yZXXISLm5ho/
ZgkeqcpmtUxutUBphfd7FQbZJcEJsWlxcmUafLQnq03fSODMfFNpc9H3EljvDx3aSRGCwS/4pPqt
r1xSgtlRBz3/6MEhpIyCiu1HSsdzf4m8mEgrdtq0QTO3TqsJ+0NaohSBqFlQCbV7THZ+Bjuj+UF1
U51AqTIF0WAF7OBKunY7VJk70XBLSn2vSfy+/tdKxtx6TM+sBakj86cDigsBZiBdkwSKUYBwiMPl
jGa0SOjR+jUou+Aej7gmx9UfAHwhaKaeHBA0z3YX1dOhu9gZ5uFaSSmcMV5ekAAU9Jp5bVd9HBPl
HJjGSgzKMiwFtsMQEfoSeKT8+Yp7KCeucdcHMJ5h64uBoyIhIpaUB6zdfhi1OEBKA9Owq6naxYoZ
goJ5z6b1jyj+ajXBeNWCMjn+7QxGxPaKQ4cYygRTl3kedqaXFv7ahsQe5gUmYSxqhTew6fKLZZf5
JK+OXu68thR1o97zG17l3Cq7m91S/ct+I7MreZ9D1ziCdlY5ZEZ5r4IkNCCwXvTTg1ab2JxV+rGy
zMJcCbN4zBnyEQ2N5V9oOY7/9r20A7XKwx0CCDqbPXfAI3k+rcy98J8VeiwkFz7fUDk4GePRae8w
G1UU34WrM8KHkGrlGNLxxp1Q9lkjBIj1pwMPnqmGXJpCJM3ZuwwOJQCHLhRPdG2nhDQZDObODK8W
ng38aa+myVO7+Q202aHfRv/Dw0GNjBNsk/2BJ4pQ9++28lzFT2MswfyeJnI0b174WlN/t5H7RWSE
wn5WkbenQ9QxaZ7IGKmltOFJmEGPW3+5NyKqV5pZKqIq7VmY+RBNLUUap3QcugzRG9QdCWpw0suT
tIRH3Luk76s/rB4y8zH7/1hD7bb49q8uSwxA3M18epsnSNSZLHpvzd/SE3a6owWg5Lh0eIIqD840
4pzTi6CuAn6HWEzfv7bk71LUfhc0SePEPvrvf5RdMXv34RGeb3LSrV20/0W+WKkRRdt8DyvOTNsL
cJ2RcvQJR1TWGCHgfrI7dnUn6G5rcbEnf+zo2FQIItOXGsfye4gW1Eoy0OHK1oAjkBbGUVDHx2FD
jwnrvyI25brQCYK1ToXo5Tp5vxOUmKkCcCVHgds6PYYT90NjI+aRLD+E/J8KHYJRZ0+qEJGRqZ2a
V+xjJ+PjJmykAZdxz8jruysGQ//9ai8L+4LaZx09WziJhgOiuzvag5U4OGq4RU+80/hfFyPD66Fr
m3S/pU/6E0uQnGtMyz413FHR0LzeNvUWO68w7fHcOBkJHAwnWxkAfxdAZ/WBR0uP8EGPub6UxlS6
4R5iwJP0HHHrIV+6HyrkLQTLsxfZh/dJ4HSz9mre8eRU2eIByZnj0O+ht890jgvKm5cmo5OkkbT7
2zmNUxN9REVmaYYMPQJrSPANfG3cd0tWcUk0TjktDiR+atDuvJiRykDNkIrjZzC3gMf9pAdLx4cH
NZLmkAxfoelHRzK+C79rZ9LGTpSm/WBeKgI6XOt2p4BAhWPUaQfGQFkIWdqxRU+9ke6TEq3R4ItG
MbgKpdJlyz6+13YCAHVvyL7hgpIkgThvqbEVhjxfW5huS3gyaGfnT4TDe18g7cFPoItMIr0VFwZ9
Z/sMaJkmd3LoS0ZLGREsJRbucP6ctMso/xHPTrBXilxRqe6NYP8vK/0txm9I50kBZkwyocnXG1OX
kUb44f3MWU7bAj09dEjUOlhM/8xUWmnZj8SSzVTAWr9LSQOnp6SaH2EbXYaZX81RSi7UIUnRMDHW
5uyXxDdytbX2t5VJx0zQRZASwvPgIxKe3zyVSGlUQ7T4Iv/nY/+e5DeM9WWcUTHTz4Q/CkUKMyh2
I7bFN2b5QDGyjZjm7Rq/sy11FgT1s8r/+F6OHyaf4rBed2jggVtWKpvrNrA+c5xxJF/4zFzl/Bzx
pgRDDM2jEMiHZuYBRnu1qRWF5me7d95YbqBjtHEUTInaNPHhR05tO+haMBfo5l0zmEGdfZtTngWU
7ACl4yr/2GpF15GTL+I/AsQ1DHfVRIT41EKwnYCdePJ3qCnkvsa0Mr3tzgXgkPUGL4JI4Sw7E9hj
rICSUpG4TZzlD4aR5RHW44Ydco2T9mQ94iv7eqety7J9NSzBqa5PzRRsb7KLSWtd58XHAHCGQNN1
3Q8lIijwZPMxPJS7+kf7FnieXAFE5YzZaKGY8oF2IWCqPEdieyvSc1Rbvwq6B2PtfSGFnveZ3nu9
glykajsNSTLJ0RjhbCy9Kt5yAd/AOlUSfxwTCEhjjDWVZAmpat1mDFweeIqrU+uVHs1m+lqCWU2S
ZYB32qj+SvbqVNaD4Dt4nfndAQzd499Oux+BnzboYhgPoMypvq9MaIl23AAyqtL0JQTCLqLL+GCA
VEUVo8ceMLMruEfwr/L0bZBb8auRUjZxvVqzWOVcWa0qnPLNJY34UoG2ZzU6wh7ldM91U8I0b7ij
UWTdQA7WgXzlhxJvPjeD5jENbavxKLCtVB9XaAGjghVbZufeIehzkKs4OJ+d5pbpJWavP0O0sxR/
0d218vVjmg1WJILZUJcxp7CepLeCTSeaUy6MfdJIidML0bjU9bXolqAibrJJeRs6pu0oEqGKexnt
+d6jALXE0M6TwAL9dgv6dnML7C9ciLKQbLSGMIdo8GQ8e1h7SYt8GNwSNqV0oOyvmfGo4uzGjN+t
WT5zPoTFg5hESHbhSJm6As/7kSFWGYVbX3SX2lrzHFZ7UyLJJa2A10V/UJtIikkdvaDPrs3dtZX/
2BkxyaPIsAL+W+WMbpAX6ZV3B1mlwBGN2U5x8BchfYAkFdTpznhrYBaFAjaUS+3MgMx3dgNTSngA
9a/VclpgISVJzQVlHYo7DYpc5ArBcrhi4L/eLVu+fyCenqMtE25gziFwOVK9QhHB0sfKo0kFT74e
OUC02FmthdwBzvVyXE9wTjCjBGVCV1mLncJsyh9gPVDmeTUaWUBVHQBX6NRa3j0mdlPJajCcASCa
aT8tZgBTzJwJojxsWPX9hzAkriekCpQ5NeTombFi8k50U/OcZPX/KbBfgbf9y441c/g014ofpNl5
hTmFmv5vFMps3elILJ2dIal0iA16ynaqLMqcECuQS30rv+ARoiNI+RDJyq8TiAvg8xL9YFtSJhek
VNdCtBC7bM7KQ2B7hQJ2bgkr3mnU9SHeyc3bCsPGABAyoijtRwnm7B0J+hwFIj6sjJIsF1Tx0XqT
YaO1o3LasuzA9X2w//5bJbACUfiG1/QuEXMerqIRGqTuFuFBBcfnnTPxwKwa01hpo8XaNSe4ZhMz
rndAOnZZE06dVEAINmPDM0C87JDlQ0HpqHirVvlhdLJkZCeqr3sQP3yP/665VtpLU983oGVUripE
iDq2oIcfZ+Kk1lYMkeITBJVxOA7e2IV3Pu4jPfpFlT07dK+9jvp41LXYOhCSxfXwqLuEvSVScQ6W
p/3VKohWD9TM3XF1sEnEK0q5JAfU5pX61qAz4U10ZmVOgKei//XTgdEsWQAbjZv8WybmPjN3pvlN
MwOeTJ3bltX/A7D0g4Kng4cJIdVNkKM4OTr2qag2Pq8ZiQWSAQlAlVUT25Q9+SrD+468V0/g669i
3o6i2Y0QOCIULC4nFuePDJR+uz+1ixigivNrarXImNqWdwSYtS3XxJ1PVQmxz+J8TgE4r3Rs5F41
2ShD6QtIVgGauxbkV/0JwMMV6wFw41OQzgMXB0YJfUYi8LTWY+SNZydGqBLZ4NyoOf96yrK4kxsn
/NQefJY9n9Pz6vdaUdKA71+RM+zs1ixQcrFa1V3JGziI//PlG9sis7X7o7HFNnNOEtN9tmNr6jmU
GxBPnOTcfiieW8gDnpJaN4pknPwG9u/UmTXsCU5zqkzQe7smnQnSblTB1zPWNmYt6q+29e+rotow
SDmMy+HAUO5WSYdneZQLSWxYglib9181nPea5bFMJx6p/OP1BAoKa8eoKENmrjbeFvlTG5sHmKl/
J46EMoCbcfMhq5mpm1VhBYzC8GZU9+Eu0JmdX7Tl8uSESDgy+I+YZPH6zv/7v03ILf/ja0Cy3IOl
w/ffLosbeYlFFpRuOy1hqdFQSetONECRj+Hb6dub7CEeSysEF4tDwDzzFiuR4VC+AoGLmGrVwsnc
xZQldt24x2FuzToBPUlAuwfXve8ALAGBtKRt12NAzW2PP9KLyFErlQ4M/sTgC/maCg7t6stQLOWX
1ZuhAu0F6L3q6/DbAECdcRrTQDtzhJiQ6AHIIpRNWy8bI3oQ416SNwQK+T8UWxhGSU11HVqH/ljd
rm2z1FlXJsnfivtYRZ8rmP6agm5G0zAdUiYICt0HGmRgFzHfyHWMx/QVj9V2som/pv7y4AsTzq/v
iv/kZ5DdfcET0rUlskI6XLiAT6fo+yQdqwNAWM5C0df6JT1j7fLwoQr2ftVwk7f8RQxCTn5XY7CL
/9s2ZyED3/NtnJxMV7LsT8dV4WxJVA0yKVKxpeZu5EG4Ch7H5qbpFj2J0GYtbGckWKnvStDUF2Se
BQF609kFjSM1yvgCDgs1seCbFAq3oTkdWHDpAEPDeLj44a47zyHIBIJuNuSkfbxgtnOlnma6yjKK
9CJaqHJcAkxGTMXB3TH2c5//qDiC9gJaD9iUSKbFcj6vOqs/IqFv5oibrLhvSDXg6e8ih82hiouV
akCPrWnjPT7j0FdIcXobeQQvDIdGkvfHLoUFMENaO6Tc4V/PjervKYVmlIBXu9vwDGrWEqyv77V3
4mwexTDhBg3KIPzahEwzB1o9+hbDXsLLFXY0vGqgR6lrO9Yo9SftcS5GVfAsmx0uS8feZs17eHdz
sR1B1fR130VobQ73qrhklVKhpSuDNxGHZ5XYy113jGcJBmtfyojhQx3Fg9g0eEd7u0T9nOWm5yug
aHI0aw+MTq2flePAP/epS7qdmSusSyJBTwOqAgLSfxzS8Qsq6bu5gyA9kzfrWoBx72SE5JCFsVYq
KAN4eqxeALfmv1/wpMQIoO42IM2EttwDGWfmz6BSygifzIIBOCtan3HE3qTnACpsobuoBklUpFRN
sN0hoOQereJ0GNeZI3d9GIPmQ7l5B+Be6AI9IG7dXbl2KKZmNgNp05nptjvXOdWFspzc5Ig/LcKJ
NDr/BxpZiErcFc0PFp/TXpATYL6pYOy9+2gP59ETl3vhTOJ8sxCjZrG61j/4qJoBa8Fdi69kjnvb
CXcjvFM08J9ZC0NahZCYFL2/z/jCno5LnRQIMWKu9BzRzWeLxT+BfbjNj6+7zUxrqqHG3uz0hpS5
2KfftFMnbuNml+5hxdgWrc/8a6ZqaEIgkpM4UKo7rjCmtnxAXye6qdd2QrNcMsGXORf09oUF4bee
pjMFIIo4eAuTuzdFNfWqQSkC+DgWOSNtY9HoQ2pmnzv+WzKSE5ARb6fy7XoxYv1G+okFKrh3hiK7
OeCcbNMbr84N27/jLl2kHQcVZvrMSTavjkqTqa0+Pw+/b2LFi6DIUbDU57xkYqOgeK10mDL258hr
s+O5MrGxzXeZwCjTH/JHzpoKrFsTtd7GE3IOrOwWzojTonnSve8P3BPNOLduZPurSeoaWG9FiEqn
eQeGeDBEKWEmGsPvMDoEL24ju6h4H2va1UB5ExPkehppGclUY8w+pcsVoSH0y/y9gMOVoC31kSDN
v8K6ro4wzjdTNmThWnxVg6l0YbbJpxa04vhE/KmwmGj0wK552TTpUx0YA7gGkSdFu9RmwA5o0Moc
9ktDEbMJ3NLNG9CAtd4N4hr1Ep9ye8aK+kiYp+Us8VBm9DWaYE6JocNSYIfOU/p5FExvOYXP/q77
0HKxHWFXVYCWJt3RN573F5CzE+ZOzZMRhEgMyqwSa53TSPYjvH+kztUY7x9Bn6ZQT8PNKjhnv2Tw
fBq15I/M572L4Umv618YTnDagYjWqBlGC5GNhDaqBW8eosoyvEmCwJ/MWbf/aVE/6XAi2jfIwoW0
WXPlTxE5+0AUh+J2O04FfuvgyjguF9B2NxcOWA4Y8GG9iqS4b4ui3I7vQ5BFqp0g8HjPqntMgu/0
T+uRazCqhz3ZHsKPkU7fyHGJPddldoHHRWP5kJSZad6Fxqiw6T8pUV3fOvHWR6qsmeD7PGAGtYn4
+E2QbqFcfxvOrRaZFHZ1w6VrdI/xH6PKmtaPNwUfrK2VZHe7yqu2qcwFluXvciG/5KX/1SjsSmdd
Iut8xhE9mI3wGqnLyI0BXrAkdAMggsdGPBWJzPleRIhtcZnndxPxtIOg89s6xo6vDR6NYZjLV4u/
qHOfQTroJGL0V2k2cGlUEN4iT3Qr4mq4bv5nij8gYzbQC7BulZnz58Qd+LJF+PCJo3YaOvSHK9yt
3bQhvOKvo1XmEkNjYgHAmePxqPkOXVvhHkL7N/jBtP9K60J7qOsR0QZzRXW1wez9PVDvE8W4LNJa
j/wreQRO7uCLXBbqqHVB2ASl6sjxDWCEspYOaDwWZAHgDUBl3glSAyM7IDcMfGDpkDw17JwDQU3M
2ZSR6HOTJy7BGCgQIDiAJjJe84sn05UfquLotO/9R3NuH3W9KqiRQvfWeRjB9sv10LqREc/I2Cym
a6OMdwaWfr+AqYQb6vTRd0TfwrQUPri5Z0eBIjzOD4NGUImJsU/f3HSTKQ72Jp6TAPyJBQnVqZ3n
4zNSZ4/DYuU5zgy5UOrOj1W/2Kl6oafHeyDQFQViATpbrM9KGcITZWJTstzmDL5k232h21dDw3Nt
xHB/m8MvEoX+tQaWttsPOws8miMc65+WbpMWX96upOteanlD5z4bkmlphDFGXaDgjgw5NtJZiBiV
63BfIPJs2rYiwZXbHwHUepxwS1EW5WRtYSc8e1896bjTTYnl+3ZzlfGohtAeYYpfVTxHeHO5M/Nd
qozxUUDQpcpNsYFcNc5jmXrDsO025CdQarb05CTCMu9taH0jqY5cf+xMmIhe7CY/7HIg1L8m+uqj
4Il9YVc4os+D4WVBnmQOB7EPQCT+ryZ84jRhrUGBwg0BBsW+PG+QDYglOvjglczIOM28RCk4JJgy
3A+u+5ct93FmfSoLOrpzUp1hF9Ogk6ysrY1+4hMiRPWMZ355jRsSH1v2TFJIzaU9m9dnwdZciu/0
eV2WFQqUkGwXacJRvpJ3yWQNFt/O7EJs4Y4+T0dVuqeXUmZqVbGLoKK0lkcKlpGFQQRNiwip4sMb
q9hVhLj8qqAXWfHC0fFRLU84sYgvYBS8ZGrB0sax/pMRq1eK0w9EVYiOI0LhZbGfnOvTf1CQVcEX
LPipBvQDUSMbzFvKPj70lWVPRlCSLf7D5x1BiQnG75PULzg++nLzrfPTjaUn1NTFVrHPNw2qx91b
m7ve8YCJB7Et2Kj+4vooNzNOi9G4MISe9OgclMqFwxt08EKS/oymmvpmLr9ITFb1pJUKDod7EbvR
roi+Ax5KcWi3VuzWeK8j/DkpPj1+02pESlAWIEQJJkUaXXmGVPii1B5uYh4tLDlMNxWHaRS4VvO2
gcPth3+wyUlP2XpBM2UImaZJiKva4PVJmdVVZWYZUtV4bsx+0vr15U/ZctDPBdARaR5KLh/z4uBw
sx8NXSr/1wez2esaz/WByvtyzSlDapmjS7QWFpeFXJfqoMXHxmtI7zEyzoauFwKCfd88+Srfdx3S
rM6wdyWnV51APG/h0VoS94+4lfFBM1LtBaQ+oHrkvWxKblNi3E9xz5b5AR6x1S2VUGOMm8fhZWCr
PuH6IUJyap/YoA8REjHh+J/tdG8fsb/AgfpJw2dCzS4qBNK9DEIBdW/F/JWO8natr60QfegxZtNG
4mG6Yocc0vc6JxnSAzTD1rwCnakP1Oj+tyuQtt/QP+QkxI7J/77/3q1h1RkkKTazC2EN807gM3Hi
u/AYXm+MGPxupMmM2to/GsEIsQXoZFDVK+Nnwt8T1tBNyW0YMaU8ElQBdi9RGyyn420wPhw06y5f
2jsThcQ84vl2zGPal2qRnENZ9+wUDJw3+4djiiVZ3eNNw0m3vNXZqpXXTziNdCsdKPxe+GUR/Fr+
YRFNEuqwzmGFMXeVMvTgUZXNdxCHJqdmu4mhaI4MLAAHSLZfxZtxPpHX1FwOu61fjbDo7teywVgd
tnu1E2o8pOmbYgeBw2bvdx5wlbsDSwva0Y9KkXSN8fe0JiLbkkow0y0DUIyfgUWnmkrBnFEWk4G0
LM/sEM7GgVCcxXRXLe1pdLVuO2sDyddybGQDUjoMZKJbzKKDsjDDKj7DwpN7opD7EPx/Ik57xvVK
08w6auS/oV0uSbEAGtq0lIxe98nJ6O9jzUxiN0ydiro8+GlgNcliLXWUIxgm+aTgve/1qRuifVct
HQRm8pJrX3QjINSqezub3ateypnxcna+iA8PXtzDmZNPBi4kphlAMYW3EIWJg43yjt0OaMMLa+dg
ApiQ21LPt0FcpyqHOqMPoOZFHbVPErtfmQ6CHtrLx9hYlA6Qknufs8P2mAUrvJLDLdQLdGjhUIT2
IXzKTHGp04ONJlJMtSi2pqQRm5BF3hSQw+vt4CbZqfSdUc/1UXpXGuXqdyW3VbC4VVNX0lia8CpH
W/fxMCpIEhwKH2aO4wTr8idHJbELN0vfghmwQ1/ADSk9OQ/ULmT/A9uqrlwkrNFJR/Wcj+IF4Pp0
EVnurUyMv6z6OSF6NH6uKGLHdL9IWWtekOxADaL2O7wS7d70G/5zQZ3HoNXZ6IhZDwn2uxxejNG6
ZshJTuQNYDNcO44P8UmlriKChaEZtEGo3xHk8Nn16n0mgAjEt1A9+RregQ/45NqQpY8y75h1UmlE
mRA8rG+u6Y/263LMiNs2PWzZDZns/yr4Pbhmq1Bt24i/GO4k36q9iva+JC8nOYjychSketAHhGHG
FLwf0bEniaC6z508rIjSjjO/1kXG06oY8smAhRFE6iaKzvwyqrkOtze+6O9FQ93Che5+tym3qO4o
X3WrsHhbXqv2+W2yR+lPwRCdOF8Lm40LHe3JcYePUehteV7AicBTAFaV5Ra3FbBCtrseX7z66CrA
PmKo8F0l7zEiNCSM8XgE6qVA7u0trYxSuNKolMxR/mrkh//Pa/9zU8kAk2zxvZ8YGB2cwK4lWpEv
dBXfF/WVA2PBG5j7NAYowdnOBG15vvnNptzPMt7nr4+AECrv7xxGv8XgkpJIWh/SJPbI674wpeSl
gFbTMAKAkfwPoRHvamEWi9tVg0OwL80eE/1TWmE0t2bbBymAZrLAEVANcWKVW0EZR702wx09aJ7L
UTJWE4AiRj3JMZUnJMkTvel1uCjHqCd5Orb134EsTgvJeXyx/gsH/NGndIduJWsQeTf3ZMVnRe6b
YHbtnfYELEYigHZ0KdsJ0g51AVOLktw/asWtYzTg9q8SJ9koys62qrARcYNE5427nJBUo1sptoHW
ocr3Am0zQEG3icajCf83l+j3wn4CtQutjPd/VUEQBjNrJvAAWnyNsnkdKgjkKVB3JL8C/Fb5TpXG
+o9wJuL4WAR0RpTxu5ynmhF/vsv/rd5+JjaVgKIADvzrQrnBq0c91hqv2vBkWkahVm9/WK3l9uez
U+JpdXhV96+XCojUh0IoLecMue2iHlPuEeIJ9IOvEVA11vO+CFQtrkpRXHjO0Wb8IsteGkDT78NO
CkDoz0wFPYULFsQyAwFXZzyvxSxGQmmB0+A/VJOMXYWMRYYUIyJ+4VSw6jwbxjnLYOcsedAYg5Al
bdiWAYhayuhugTSQiZsJz2QqA+rLNx/4do1tFTQVkJd96dYtqzixUkL6ChVLYk0HkMhe4xeX2MLF
rRf20ufelYlwz6iku3Z8hEWPOBZ56m4Gmo2P3mSz5LjCxqzv9CxpFA+jLGeykkO0bwQcE9CN2J30
lI064dfJBhSeusLLZBJ3XhN61PIFoo7JazGB9fupZRI9+U5kSDp6bLxwLdFsDwJRWhiZueaSQPKM
t7hTKZ5V6w/XW7D2V0gyaNr52HIwf4qs8qGY0KcE1kfo/DGgKZTEmf9icIUFVDsqp+bprtQLZAXz
TpvOAcqKA3i7/4irOB1qLJ3kGh0g0MvRmr57kXd/s4dHuScK/NZECGNyvvmg/ZVX7OQSW20YRkvG
wXVPh709p3lV205pSB2U75561iAyX19jRaXlPZkqGtvefVDiejjYdTTKLjvtqCOXFNnNk4wMjjvi
gpB/yctjJxg7tqHwICmncLvbSGEYfGmrfjMH+VZH1AttbjWbQ33/EPVovVKuOywfZ51XzVShwzkM
Z8OvWPrN809pwwwxEM59nEWLmZMVslIOfRM2Gof5TVfHDaOx4T33yPw5LaKWoEMQHUQEqnnj03G4
Ys3Mt2nBfWCIMCk7VtWbbP6VkWRvv8PvpgHrGO1egK0fp78w7beBf0m90bbvpZd2UoDHf8uHsUOf
rTgwrOTbq29Jq5VfEJvTCaA98bJcHCvT7xw3XXPPDmJ3hcXcrMQMN24T+YWsyZBSoeaO5Thmm8Ya
UH+XkcEh8wRQ8rJa8ET17nTcSDQAPfGEZUPnMWSVPNYuGPC8Rr8xmt/lslxMHn++6mF7QUxu7tPm
+SWwj22fqY+f8L6ePOuP8rI7XtqgkngvO/4lbw+txYso+Tv86V7mGGpDxzjWsOkNXBi+ghYl+WLi
SdzQlLa/pWWZQ1j2lDXq2jJw6Ld1ewxTZ5TX2eLWMksxahMJfZhr3Dm6Ykgh79gyweF/o6ZyuGIY
ownxkEpIwtaOiROslK3PSMLKhH/mNtRSeo5z5pWxLqFWRJeddFxJFk1E8BtrQcsPr4bNg3au/uYK
z5wT83nVMF3bW4yt+O8IJRzqfGbvzzaTuWxZHfznJLhmTMkO4s0eumjYTROo0mbP/5fdTQyMOOnL
0yIBvw4gLLRid9gdVFQwWAUtnVhPYqmHoVVj/Ax99pIcquPrLHE+S20N+WyhulUYMrRFm7xooRLw
VFc8lYH2d+e37MjPZ0a/r0WlFj9RaZewhL8rWhrcsxjGsvzNV2s990BJ6dAqUv5/BXXXpq0uPP8r
saGp+t3ZvUCkrr/aKlC70cKlv62I43sd2qYogjhFHThyg/qbi1QvsncUrvFOom4I3CWzfJSPWF4O
PFlCKmPA5EylYQ+60wkta+sbqsKMwJYgc8aa89rhKwKcBbjNHKuVtIIm6oAzzIodOg8jv1Zu78g9
BFUuKxpoJoPiDfxfaskFACmF10c2vMl1kamOxgx1lPFbxl3a07XC7x8vrkpoEv5yZm0+4ys/CwzM
R51demSiJftGZHdrxUZPg8alAE1UpWfvUleBcu0mcD0RyShbldEifTxbj5ZC2MA99qPCpp4iLJK1
uXzYPf2teAKr9gUqfzJssLwwjylaFvATdqbW9fw8W+alhIodbOXZn2Zjp9pNZXqOSgMY0WXgYz1U
kGcYGYh4nU69qZ0g2vw6eJsev5TiNVuxF+Hk6zVFh/7bWp+ZcvmaTBarMQ05/wexcF84zzwD0PW4
bCeGyo9foVtMFvvSVlLki4Or9cg3NfR9/SwNOaVWakBCw+oNdRR/JZ40BrBkpFhCRGa+YrRAjEzW
iOLoMVmu8Lu4OAhHLOuHf6Non45sg9GWYtOZijbAVrRpTaYomXQrK4U42NrEuag4ZRQ1Od3aBAXp
WoOG0YqZoPSCiKVBru8PY6U50wU+7xkNj8igbuzKH7EeijS1vZCoGeXnXiqvqltCZegoTranpncK
hcrxf2lTBF34zAgERVoLlwa6vBWBi/mGCgQZBHuirtIZAPjABUI4yrSBG89XrSbgCL5mxwj88eAY
Ws2dHb9vNMpCA/Wlo8yH4/fQHdHhD7+I/8wDHgw7oMg6iVZL/DkZulOKo15FAMfzFGAq2CKe0Hdj
KY3fQ8IKOZk6jzDCYfI+eSM/7MQPyJj94VvPX3FUpEEkeS38cw7VumbKZuLa1OxIrAewTohODOqn
Uk0lT2Nvos9zTEqEuWag01VXEL+TyJ5uy44RoO1xwbb+7fq11SJvlGO/1FRxO5uXHYnWyfoEpELn
k01LpgOgiThX566IT+RLord5KGKE7XO/MBmGmQCrGtuwDxO2VLLOGEkBp5gHFQid3CuzG8BY+8G0
UuD3WLAoJyx/gSGOIwrQkI2z+wtaMD/+W3q9XSyRek0IwCrhIAajY7WFJCfABk9c8tjmp0GnhzGt
fasbAh23oApRdvIb+CT6xzPqlvtneI4KINbO/Mdlaarhpt7MUoy7hmuAM3CLQ2o7/NezzX3ldivN
c8uZjDZ5g0A+K5g4D898P9e8qQ99s9Braj46PtSUJ7d4ODR3d5Dc9BJcgf5mEp1rmZxcC2l+kv6j
RzId23zrmp8tqchLdptA5qWl9vwK3hNIOeyKL+pE1MqRIDwpPju/colSjUTbhXJWu+CCDzDRqA2A
Vda1mFTlSDqW5+MaWk1kcBfZjYHLOqZroZYfuGnDX339ewEhPU5K+/OYGt0oeX3WQJdMGcic05v2
wKh27+O0xDOPEmqUPaV4wYD46c4akioMA/p/FrBW8fmX5c+onvwVsIM7G269YNtcZKteh/BQAIni
+UsuClCyuykedU4q8WufGz0AEDSsIz2Uc4RgPfUP9pxcznGifwtFSn7Vgirf4cnURvsuwuNyBMX5
5D53dEGyz6AenwdzkPe9X8Zn7m6ibb/n8k7egKCBqtKaY83Ib+hf7CYEy97HZTKwuhO25+tyqppJ
hjg6mIFS4wVTa/CvvUf3jMfbXGT3BukyFIL/FW/cI9cUezec3A+F6kRBSeUnTnhhFHxQ9TbOj70C
U9a1/FfF6MzJDtvVPiNZy75nP+qFddFl7xRbpkTptyccDtTF09lIxhaNkLvCR5F169Zb85e7vBvU
4Hbyv04Hm3wYaxW9tfXPV3PLGjbGbHqZoqrROcrz8Fbcq6x2LDKxdM/2muMo+DmoEMYSlN8n3K/c
e4qIyWkhMr6wPT/himYkJbW2uB0qsN/mMg0ZfVxfzkAxyb3LFpecv5DH1LoeiCgUGkhWXoLr8VyW
bDfcuh2t9Gyjj8K1s9XinWeW3+C3rW+KjMb2Ig3BE0vp0a0AELM5DuR1EAz34KLYjEkYhEXx4F+A
eeaY0pURIzO0CJvg/+3rdhgCooAUD8768hn5+8BjmhZxY3UWsHWQQEMhDcQcIHIl0iaMmRvmE1/+
w31Ww3HaAiTDK/clWLwqyVfQmItCOU/O48LEcIxp5mMaSovfgmlKToPpgDEPKXT4AV5g2aYvUS8K
SQyw9/glim8ecOwKcje6I+qpfABC/cw1jwsFdUr4z+6Rg6/njJJOPGNAXwHgjTkYCk+kCsc7cfEr
0y6FD9xlM0aRBWTwBgj0ErGrr2xBVChr5sHMH1abptHwFuMZ0GvkK0wN2eWAun1FA6ePKEfBhKPh
UFAPxmQssZsM/fZa5EH1XAmJMJY20PMLVBvujOhu8nlZVc/xHnkVqT9O4HELvwIEjV3JzrA0Gs1X
M0UZBYuOLKFx82Nyxb8KL/X9Y96W2oWq79N3ToqecJd7z/eVjCGHlDZg2ia7b3u6DAIiYQHl8RVb
ej9lt5Uu/YZfLrjIWzuiCWanUDDP9fXyhmoCFDUGQva12Ysr05riTtBCnnr6pzPG5OzyLRdz9uNi
j8/UobGFL+RlPUjUTGwjsylrfmOLLUL1h/6BGBxgv5NXoRcqTTLX+LtcKSqGqXa7P+t7qP3YLe3H
XXppwt/2N8KLwnPoi8Fd0IpjSo1ROPSMyuRa0K7KOFsaZ2Kal8RBx751VZ004CUx+EYD49K0MLaP
Jyq85zBMdSFsg/HQm/iYzon0O9i4UT6DbqnF68nfKEO5ljmeCNmiV+Ot20hPRijRF97F/1TavGOZ
/U+KCw0hVcyIIHb2ZLSeT0aDPYsopgSKKPI+FUvBVzup72Gy9LIZFYAl0y3CFhHDj9c+nI93Vh4O
3V5SPOP5w0kK/9aCvw2ZN11ddZznB/yCNdtfTpIE+piATudymv6DQWReXgk9cL7y/5uQZWzinHzf
CeEMznsPRFYqEKy0/8zd/dHRo7DfckiqSw3KjARtm1jpr8bU+mf93XI3qwSwAmTWDLSCEe77uiZW
aIp0CHB+sBDMqi54HR1rt2WWMTFi4dUM4SI8Q86Y5L0ERoJahr75wKAj7tNnhMuqUuYveZ3MhFZJ
RLwx0Py7U4Sakp45q9HcxGn9tqv6kXlExA+FI/MeliaVlZsVj8YCGxONtobrt6+wF9eQazUKDWlg
kETzqaRWurVMm6ZNeU8JVg6QvFCTaJT5iR8/BnnwAFRR1+uO2/EYfp0lsmFmsSs5IL9lxBY8spsh
l/o/8Hli7VJEa8bDT1UR3F/q8+mdHHUjDEfJR6VXZXx3X1uPzurmxRIxyzvmdVaDRO2jV1JgoYA5
bA+AC6uviD5j2VoBpu3f6iAAQI6laTrS2qrCyXQ8bx72i7h02oYKJ2RbqeyWUM/1AlCHuvZ1K+0v
1BAW95xEbe/nbvMSnXGnN8ePjL/BvGms1Ohvyr2XcNOIlmH9wpoefxMpKKSO3jA7ySjXqLijDzve
3ecQCjwb98MZ1FT1MkkatCyRWL+1T5bQJpYVNrEA/UmNTXRtXsbk/VQyQaF0zLMjN7yv8C7m2ilb
sVNPdHncSf7KNSENn9G91VIvsqHrYKVBctahCQ5gijXoOXIZZNqIkyKRFWpugVYkGYbbM+RSzSnD
W+dg1GsYAdI9RbRUkqioAXsgbGkvfa+pFCYKghUw2bkHxdbdKx9K4N85Bp5lns21k/ZM8VTlkGLd
h3DFxapw1rlnIoz9968YWD1UOwtaOJtMrpKlFRzr4LMJm4px6NOICnyBbM1YPyvAHFTz2M2v8EjG
2Ya53wskOprdV1fHAE5f9U5GcleE+dyCn7455DYRyZ6hMmBHHtXsndZTfpDIuIra8NJGmLd+LqLJ
133F1KRlLJMipJg0W31K3vrzSCClRTfmBlx1f6Fi+iCn5axV94o7rwi+LHGfkulvkt5PSrayiD92
b23U7akaxRirqGrp5gABYm12n7lHsmoI2mazkKMw1Df2R9kJUKZ2dNiSjZZUSyWpC/eA1IIMQiM5
y4ygyyZAIsVkSRqlpj5/j3hP41HNGb2sBBr7S45yKdca2fJ/7yjrEgOQm34347wsIlHmQqsFpgdf
dZfpAKLJgQcdEL2LHzOXhXQT1AN7HfharApYPfhHBuf7L95Z0Yf0VE9UDNBxw4CyBUXJaxkFwc13
qvSIjrV1Q3KbcAV14p95EQRQIVbI7UxmXKzOanEXllwK35/4m07lgsPeswqvTOzHiVB7OtkSfjZp
yusOTBtjd9h/aF7H7qtOd+ZWPKHjn+YQNAwD+dHNP69SyX3tXxRT6Qbix9LjMAKAxtPETIfgg0y+
EihcPT3t8NWBvuRr1fQco6OxlxBcpxFTui9PdyHI/bCaI1D8CE/hmTXfg/KgKir6GH4jau3PrNHR
s8zPOvbwZAhyu9tYQU0KSLtTYUxOQKYEPIzKe5WE2/TsuyB3Rlu5YaDoHxpiAY3qHEmoZB1MQSXD
/uYBTAHngu2ra6XWtOdfdTXx7hiAOJ+fzMvL6q1iYRGKhYuGQ0WsOegjsQZazZynv0Lbab91/1lV
Qjcft1+l0JUIvE/yKvxRcN0cVZyDBoz/Kbi6MH9yw/TG3+suouchzyxwf1Qcp4nES5DTc7s/FVqo
6GlNQUDpltOKsKEB1n4IgV1Wf1tNoZxfMjC/syukfwdlnqCWqMO7NfInLDwS6EFD/SztVSzramTu
jlgzaQdhfz5DDFHtn9gurKFr8CAhzxFB/1bSG75RMgLjTndW1mWtX1vjj5c4y2rxZDPoRS8sjL2d
6vUMs/atvgCNb5++n4IC7KdzKPHmxZ6uZ8fFNr51uuCEIOTM/7PUQBeaJ1lu7P8j+iz5llhno0c7
6uFdC7MQcplVDevMNTrETdyenufavPUVA/ceKuUeSDbX4GBtPGspcA/agWX9GzbK3KtI6jpCg/Cb
4s+ROlzVhXmxwgkRC8h9LiWIkedgjnlw338Nhbdfo5nbkX9lrEkThTDhIByMVYTN4gnGXWA7TWlj
dEDeCg/GSv0n8+xCDj7L8wbw1BzfZNxpnrBttfErbxR17RNzJlLif+PaPP6kQWTO0aqAeH0Kvz2I
O2je63PSImspEtLV5vHAHUWE8MhbQBQ3D3XinCzG+VggDtewBJlFv4MDr7Vm2+ffUx7KrieNVuqJ
Z6upFQBHlS3zqNXbPeZPZlvDjpI7tCTESMHZxg9/zSOr/MQwnxuj8DhGY+HRpiRiJbhepXfK2xPd
utAz83qZECwBmPLzew5/LbyWITR6P73j/UrQvoNYg84BYCEWJrWRFv9HrgCtjltOHmcLjajqXHzC
O8v27IAYokIwiHBwCcBcKMecCg48oBb7Pp4A1nEWOFRcUFiVWnMysUqHlVt8RGliwykTBsv8jGoC
XiSL+H9l2ScIScttCiqtRUrg7Tq/PP3D2bNevvKGBKIZGQ0xqJMlIIJq+XlUgYbMnOB3AOFhbcMa
CnCNng52RCmA8G8K9OpNm8WKuWZtdj1a0Q0ysrtRcx+znLBxH4d0l6gHHSSowK2yzfUkVBvQqOw2
eKhEbUYq5weUASCa7GaEDXIqrCa0eSJjKf7Gm06NnzjFUqV/CzRpLerHR+VqCTztdJakE9GD74TO
o4+X4mZIFsEbAMOAt7nppYuFrxgm+bxRVno+xaW5V9JfQMmP5fnz6qLGvMYayfBC0hgDUEjrmap4
SAobMHl/Rmiva5VF5oHB/aIfVUMP8mKsp9wBMd4nEOoEqEssVwa/4hdHA6TNisqs4fRrhVR7RvqI
oQkNxhF2vRE7g9Y15NVnvZ/lQsUkAANmqGlh6wi1xhuEHpHBfEQPEk/W5wYVMvYZgrVja1wVotN7
r0RCJ1Pqk43DtLdsZMLEFj82LsVRSEnutmqO52Rh2sW1wB79CXHDpl4yPIXw/61Fz5P1pC4f1P4w
76lY/FAHKgfQn3mvFr7B89cnTxnQ+tRNs88aqEluILBY5Ek9bjjrR1+yq1BZEISYewzlNXK3884I
lleazy6OlcxCXTlj0QiaCGcTswNM8WF0fyo8TR7C/YlI9QteGLnS1ZaNg4A33WTg5AegnacyjuSI
kwIqlAgVOM9CzfXyYNfwsu8uudsVSv6Wa+0rsSyaCZoKyIBOzHky1yGYpw9qnLyx5SXWJntxbyeq
4wlpZpbOvsbD+ju5n0vmji4dclgT4JiJMx1jO0kZx6RICgpMnIM7eQCC1SClq79SfvYppavGnkzf
xk+m4T5udCfRunLpdovmFj+bS54huk8aMnGdBYPG8FZTjgNnxXLaFdjhINfIjC9JrApXXRW7QaJo
cY/oWupIeq/0a+S0a8eTJFB0sUhV0anjtn2ixGQy68HRE5jGU3yFmC76A/VSqsv2QhTNloS4UgB3
63rReGV6mHkivbjRoJ4Jw6ZcavGHEKLz46FEsEcqTSSeTmmzxJMrnuqwx4nPLdBqLy6sWETqh0G1
CrlE+mUqgBz8Kaw6GPCd9PpfOaQSHbhOF3LzW7ClH6dPrgHjcVEV6Gw/J0x9LSWyV/9jCHZu31rh
N1sfhBuhfUPYEvesFOeulwQ5jizC9qox0bQX5PgiYAAGzL4auEXL6GCWbTWTCXTnPlAw8zTTT7NR
VMlcDYy6EfV5iA6KmKfncu6DhY5qZa8PDQS/Br87mBwl54EipiEHSgx2VpDkulK+AJTjGHrJKvPj
jWtuEoXAk7ltXvF5YS8tawCS7ZaPW9FpuibjRN96NWeeCPw9WKKe6NLlS3+wRR6sp/7XQe3wkZCB
so8VkBvdzsIOFk8sIA0jVC20ZZE6YevHFK4MZyrlhrIm+0pVOmMkKeLk5jIynUQwajZuv3BYAki/
eMe7mii1A33y+nANkX1ud9xZrGGN82AxG0bO2JBx/spaaEyMfEmZVFsfoPcgx06hVBHvNMDQqISq
dAoMNlliEDkGx/Cdjwmj0MOGop2eZsJBo/PfngrK29dDyaNmYh+3qESfmu+7x17c4DzQp3oMYItf
oLueJL/5V2qPS52cOlyGt1wB+iIKReQ2+gWLSJd/3NCvVi0xohDVJ3u/hXoNRw7bH/e/fKEKiJeS
lACX0FyeYvn5/928y/2KvB16IRC1WoWKGuZo9piuHaYYjXNHmYW03sCx+JWzyb/qef2Ls6iyILsi
WhA0Enf2h7FaMRzpNwYpampLKo70pTfTjU7AJFYXVrwz15f/on0zFlOQ1W/zIZgzsNmk+rjotJmQ
m45Xome1r413JX0CCJS/pQvq4xJpDDQT0X27TBoZIAEl9ayKKiKYBSRODeXn8RUF9VbKxvRXjkHI
cDspFW/imrsP27HN3FZdMKxQOkLaQnz9w6XMAneEqBGZSHHVKA1/LPcOlsE8c1YjBZDMNUI0WkXv
oKlTFm2D3D+LZUFkalrLojb3bwUEKWJ4IcgOXt8kzkxK0GCUiveG63QB6ww3jHH7jicVmORchJbi
hDYivLf+ZKfbjTdqj4DNLmUa7rJsoarLwf46VHFo0CtyM4dv/d8Jn5Ur7Lgt9oWl69HveZpA66qn
2CDBV7vN7p2h6kwBcqQEQR8LeGOYOJb6YXZamJaP5mX2iykue+felAuA3eD//yDMAZcSiRUu+EyV
+0cMJZRYQDD9UIYd7LKzLaMcboh9R3lL2u+x/QqgFluOQ3anSnoPgZTh+uiSoHK00pNqiwn2S6so
deBLCQPkrZ/d66q2bhFt0XgQ0kDxpH7WIKBInmEWLw6yLSbiaM1QBrzXgfEMlSEaXGKKe/JTVUln
Jq82jCxGh1FUoLpZCnGyEnojhE+opYOtcfyiXbl/SF9Ng3RbSdLNF11HkaSBdvmsD2Wy0kYmi6VM
DUWnj8htXKlri7EY77f6Qeb72T4xGKmrD34wW3YcmPxBVj2GZIqOE8b7rOzLN/qZvLBpfvQ+Z1qH
I2sLFpG0IcAg0AR5svffbj8UfAfpOD2v39HFglo9D3PWKULaRxf4+8k9WxHhwEluqHAwXysXm+AA
4HglE61LhZD0BFFyjv/KFnsEQRF1yEbqqVA5MCYXpSI0ooJbovIv0xYCJU4ZxceTwwUzN2vthTq7
ZAC9seblNtcEBaaxraS6ooELwejMCIMsHfUrSFKZdGA0+j+/bvXUy6EY6B95lA1kvEyXMg/1tHlF
IK7qQgsJA0e4JqNnqYzLq4m82nq9JaRxDvv47yPfbbUStueYa7+XgoJ5z0PHsI3e0nSNxzvvfjnx
rpWZ1ZO4Nv7/ovPvAzLbbnNLzQBqyJ7nJDnkXkP5gPclr4uRK642ieGgQqKu8v+yyIa2TTgiDZDB
6R+iR+qcYOIyVRGjglWj33PkurMlveOSrzQSmukdkn7tAcqNV3r1vlxsuSm82AiKjEqSNEECnWx3
g0wcmqrSRu+EBc+6414NeiF9nhaRVUjVwjdoA4lPv996Kdq4Sszj+nLn2H2F6adnpcUPXYq+IqoW
jPsQbVwQKBn6tIowjksGbWJu2Av4naGFqoJNvwLX0iFjh2+do5kXQm4agWG3o1cuvDZ3NN9TaA+E
Ik1GgDLWkn40Ql+kd46RKPHpzLeC+yz7r/X0p0/mN2ae/uRRoGlTQXceahffOQiDmFrKfhuGhz3I
Oi79S3sAlKQ77/PDdBluxQ6Y1ovuXgahoaXdLONxYbKZrI2Ym4URUmONho4nZHG9f4W7gd8gZjkp
k+t6YrgT4d7KVJbIIuhAU1NHO1H56xgcS+Wero9iqHMCDra1bKknb0p+szt3YYlnTOKS1M6Xru50
dTEqH7C3bXdOEdpW6COCWV8ranikO3xfVzRH824eMQrvrUQAxClC2mwA0v3qIPocZbf0+y4Ya26g
WE5hXx6BAI3KABLUqWzBXaU/F1dynrEJA3RyLZQdyzTu5f4VuWn2K85k4CM+j/Cc8WLmcNJZWxhI
eZGlj5QB+GhVg/R4F10ceh/Y2DiRkRxvKBJ9BOEL8l2/dXKThRnfQZZH70IDW3x2Bq2nxoY0jIwz
TF2mbRFj+KO8jDn4e8bGVKd7pkRAp7HF0tcqOxlEyYwtPqEmAvX1Qz8gJOrixgvqk98ST+i2GbDO
dT9oYGcQZS/gHN+zb1UeSmktnrSZ/128I9dX83mckvNP+wM4pDG5V41ZQtpesD1v1vFvlu7ZfGYb
bDo6+bsFtAniLNJ3NQRQ3ugnI4zVauVaHgU6nhJSrrCOmtSreFVwEE2TUSiiDCTdGQQPBtLv9Edx
rSW3fm5x/2GkHGwfgglgMWNgG8ZPP2dzL7CcbLaxiHUINJ/ItqtBO2NcbBnBmOsng6X1zDaRTDGp
UmQHbqraCTR5lqZ1kWxln9XGbQ9ciZWIV+fPS9fvqmbrP/MtRTdoR1JyaHdGDxTlznPNHtZgnNgO
1mMeimXBWsf7YKg9a9rn2oHx54fyzqrnm8yfEYRAbUhG7YHzBlsvbruEU6NDpk8xaQTseC21JqeL
MKuMsnnsNhSgk1LLind0ahflwDyYg6Ip/P/n5vE/C1SUjZFNVXSw2xqhYsLy7Tp2w+ZlgvVaLXkJ
DKwNq2timw9sff2DJYRKkVwFB5AOrSg0xCKzhwEuQS+BwIRaA0NozPVAwD7zT+wCg8UAMPHPRb0Z
3Gh51/kzvLSiOQiy/rLrAcsAR+lXa4OmVoG1JF9S6ImsW12ivk0ZJDSZ/pQPiJI79rZGn0v/odMa
0Yo2GD9tfkNMUERXQ17fCMYPpMKmzkUuYlv2ghAu4wmoCLET4iMhS8kGu7UFV1AHgsPsCfP3fVcn
blJcNCT759hmctss4CL3f+qbv5d3Q1w2f1nko6vWeq6y65B1+xJH2gJfbZ3dnwDMu/maGPI9H637
TqyAddvsHoH301qHuEZh3d1UEKvaN4PkjiK1yvfucgrv9oLX9KwhjKBdw/guyVcaWAv5LOZFOM6p
6l3aiz/BlQBhT6QGgThTg2QPkxYVCefp+3koPf3TV1B1PbLUQVJdRQ2715lTWTEHQPRzv80E+4wL
60YK6NZJi8qwcogfPgXORu8ahQs0Q4a0/QAPskMr/jb68fjduj4v3VvADsMTnhAPfbH23lB7cSxM
ir2stRpNTsTM9drq8LieHcIFbx+e10Fs4q3Ow9ohnQrEOY4OKWJ5RSemNT4l6Brzq55HJdxOQUqp
4IuDDDv4s15oyCtIJm3n61tD9wyFKmoCZnyEkEdKucN3Lc05+Yvj48vCrD4pf4vEHX4mMt0YNnV+
99+ZLMaAJhUESUbJOETRHKt/a2u9D1TJqGSXMXr5k4m2Rg7iV7P5klW2d5tydr4uLZqqkHDuMgQy
sKrfkQ6J04RWXtQb8yX+66jK9xf3PQX/jbQA0S2NHpVATWOOqMffuQilSuVnJyt1k5meOyeqii9C
PO9apAxURanIEFydGuPlugJsi9aWg0sKJqOvBIM6ZKHzMGu0NOPtDcNuM7za2GxzxCNhuBLnZ8UR
facm6D94j/EB/Ubh3SQI229fk3gda4TkK4AugDnj5mw8b5yqATRUWfna7RrGWhFCHsEHsquDe1bV
uaWmj2habbXKrMmIC73kZ9blzMwP5RE72FjAH5UnloTgL9jBQeyzirL+CJU0PghzDDsE6a0Ris9C
bkQXoZPGw8aiF/fZwJCnlTFYrnTvDl51QFc6Ojd9tGUs3DsDQwx4/FxrfwoeQo8c4TG9ZT07LVmB
GwYm39wDLoFUvjmUn+mhV7cLsovgFZQTv0YHiYlI4SO27mZd+1f/+GIep8uHHId6TOQwPTljlARZ
EAVzsoC/9ZxLJfblAEoSmQZC2DmybADvcuzEJ55sBjGT0HWBgfiCYaZ0WXexK9gHGpmyHQ4uJcGE
WDhW0acSDjpsNhHp1UuTq8CyxuVAh0OB73Tj9yovH5k9tD1SPOysmnd9hCS5J+RtUSKhQkx7Fj2W
laZtB1d7xzkafQB0mRhFihx/rrG3vbygpgqp/gF11HSs0nGNU0SNZK77y5s6iRkkl0fMnBT/tOnF
yxYydxMxvXoRuPVSjmT9mvAKxEkQLxtiLnhMDzHlp2I2U00vSEUF+7VCzGl4K69qvVBTloCRlUtH
MxacyAJHk6urL3AhkvS5pC6oYfmQRNZZc82mFTevA9fabzlOLxsPz3+nQuilBcKg5ZK/+VwtTjAt
fbMcCJ4J6UgZ6teJp/pK8mm+PnwjyhpPjnF1Eb8pbfgzE2cTKVirF8f7ddd2gsYNdZvzDMUagrKc
yYFYw06bU/M45XmlyVIPCyhgZ9cxDR5L5NMQ4Po8KxA5XKx25RWbjjEqWdxKn5q74Zsu/sWXA7Dq
RVN+djHYFIkGAvrVQxqfsHXTTVY8KBLKk/+b4HJ8PkFSs9li/2/2LjKy+8qRoB+wv30yUxi9TV4m
FFoyCKLhtVkBp6VIPMLr4XKMKVWT6tookXSdANEPRc2EJsecQVG15UmTcnJBPGm3Kd4970qDAiqZ
6Z3wRT6qi527EsdJ0mJZ49rw7rIDS5+JHXs17BZZfueJ+KnXwl8c4WYXJXdgLcfeqsiZNA8XBADE
lcxtsuKgBkywXBBE6kOL9yepsFJ1zx7h+zgOpC1Y7cYqkaSJ1K/NLU/jLrGR4ZWrMF/RLgFSzL9n
uVFn0AR8Ho0BCWpTU7ggu2uZfPwKt+yXMfXRm7209ugLVFMqQLaeie/iWPUHVyGmlSRmZYftVm8B
T4bRuBOAXL2l2f3j3fYIXZaFQIUR1Przty7jerY/k1+zEK07OMT159XFHzCwgp0I9nJMtOMlaj6y
1K45m0SGcB4KHJqz30D4BiDm04waycc6Y/9O7/cstt2h4FK29T1lmVNqz00rHR9JhGpZCPaKnzQd
o2I1esgv8WxxuZD1M9TVBP2V4GSbWsDC8IYF7nGSJr8lhX/x8g//XcoCvCD2hW1vSedAlPWe0Tqz
69K3wIiUWA+Uv2cFeIFMvvr1/rO+E1gQVIA6TszqCqJjtW4KQgLXCQjsGh85AYIoa4iY5GCj3vIY
ouAOcKu/2WPt2oHbke2HoDLlPStLbIMDYFqbQ/iINI2g27KksICfc/SV2cUEyyh7HnJwBN3kvY6L
hXCnCy4w3YrBgqREOKfZ2OxD0qsth4mrThce4cp1kIhZcI9o8oKLewlJminQPviJFA3ECWHBgjQ3
k7ZvxXH4S/y/MNhJ/+JMbRa9Do8bHI7l+x0uGedCaVbI3dXjbwfJkIBQEZFsBJ7w3jyBm6A1/cfZ
yiv23p54z/ZZXS0Hs/C/86R136nRtM632G4GE5jlwZpU1RsMRamo6eWOWP/9Fxk8t6VqrxACHnpE
gRuPU/984Fz1tTOaljBh54kOKVi5AmZ6XxdSxsNejvLxsagtksAVi0vpf/RnNIuD8tHA5xpGBwhW
q2mwUGAuVPiz6cxhRN/TZSUJU8/GRLOuqibZuHd+lWoENK13Kd+qEpXEgkbaivkw9PVFqXNkL6O3
Fi4yV4lo0/EFIgFHdlQS/l+uDTuzXT6foNmV4txws02JsttrLYJmyddaMXSJ+pky1G5lkqkA7ojG
36fJ9tXHXn6l7NqaJ/Sm1Y0BjuzRuC+bzzAehiCG3VUiIXdpSfHxkgpJ97QKp2znm4iERT0CnuAw
JhC+ZvFHCQSmMSC3K3eSSLw1hIic96UyihcgpO28J9YCZuTR5r0Jg7wQbpvW9Sj+EDeg9RLalJht
Q1cP7LmpjIacDiX/2/y/35b/mE6qDgROfV3nEeQyVQjfm7Pq+576r8arm8g9QqvsLZUbq/Ol7C2m
9O3Y3aEtA+iMV74CRuXiwKML0hY3GEjOTL7PEp2z6dzZdIDsD+aTR9d8EG6Ft1dsVFyvFjXN1lzf
zevUrPGgrMsQ6AFbRTpEaqARxKvyAqEUVNpW99mWbS4pnv+H1VzSkz5+KZMBtxT5ikP055Fyw3hg
KddVWi9C1hVtPZO/eA1xQrjQaWdHIUKxQ3Uoz0BADvN29KHeMzmzqzGeKquHZNoweF0CB/5/MDOy
TVl3ZtUEuKBBYNhwFXshaKVSL+Vf4Kdz4IOifw2e6hXqMIulo5m0a9u0ltAzHkMIlxH7ovzbR9sQ
kRWwDh2HcLDu/1SD4bfB522I5bzmitwQxnsTfagszv7F/o5hgtkcjVjO78EUmTc8mqVNKX0SUlTP
8q7IwHEUPHHLBh0wiUWdSCs9tLYZClhc8UvV5GoPonPKKIXotrlefrxKwFC/S2/oN9rpC2ifJZqU
482O8TB2ET77N6LKtH8JYAghJDiqaBUSv7JLog8c5jo2RymOBWizoP2xrhNNDRTmmOL4uHz9d3kK
K9WNS3nbISQPDXYe70SovL+Vbplk5RexBtgx2BOSYBdBE5nnOo4kY81YO/iIt+/A7pA9Lvos4hLt
eaafEpRYhw31AuetMt/yD+A0Ndih0isLJ45ZAUDBa1i/Rxb1i4TAVt2SzdXmV6Me5gly5EDufDrF
1R6UXYNtAOD/9SPx9WpzxTxlvVb0pzbDbK9S5DqQbiIRwdk8kynLSfsS65y++kV9atjAAO4aQXGp
seciMD9vl0L4quJYxjI+m/jzcnlqj/YUSxfrPvmKpCYsptXIKD4jZmxXe607Ib0vBGlvutEExgoV
OS7VfOuiahlLkzAfA21nYxyUbkTLeqUO/qVjoe13gLzt5nwEssRdOOJBxTUntQEu8gJ++WO0ZqeR
VcjC/IObRVagfSWVHDwFlQmZByg43bWaM7XgAPgkJd1+r1SL4Yb20DhrH8vb5YT1OBhBtAhRhqga
Wz+5r7n4P720mICGDxJ4RC0faJDmp8L9VyKmkoQiluRIojFUasz8YYgwqc7DS54bhqZXAaRe9yra
o+s0hNAxjPApCHVW7XJ2hpvk5hKItFkGgT2pqJzheZWHGzIPUOQJ16+d6y5ngH+RjcjTCeV7MTi2
WaOuqSWiC5h6L5ob5eULrHlXJ5kPQyEj+m3IhkNAtLTEI6/ZQPskpR1lK7w6zCml7bKSOGP49rvd
mF1tRtnSjKcadREXt3qYx3Mv3LSMlQJgwFpJUpz+2zjBlfI6wHzusqX0tC9tewHckOAzFeiTe3Ge
u7EpjXx2I5wh6BWiRxEbuGEoTfpKbMOl8NNOSOvl1ySMHyjcVWmmU8XkPpqGegLv4ytTfPWYjFmb
Xetkxe5SSucFcviWt6dM77mnTv9BA2gSYHP+9riH61uzb/fvt/51vvkZZeDQfjcuSUYxBgydo7RA
AzDtA7HiCMIkF7AZxoe6EhxGOlOqhTNGR8u0myOLt1sOzCxN1hJ3Wc1UoSzA4KOLF1HyuG90yTzx
ATPXS4uSpCLeJ+XJyuB8Le5PnyTsHL3bXPzhAPJ7MvXv2z1Pi9ZDprVTOI02dhhe/wNVdUL4e+9j
3/aNirAR6RoYG+Nx6WNTrWQ/G0cgpoeT6SwA2pap1E+Z58CmSEKVz+Gq8u7YbUiorZTlzi/uyEE6
79Hk7cKICSynaWNvuPepwSk18Ye5sZYMgnQtaaV91XfJZyfGJZ4ivfyL7pMktNy9OWOKlQuZNurw
zxNEpxeyQJ3Oenf0EDKZT4ChUGpekDi5KhGMYt6VHar+ZV950uD1bU+ZTaWYJ0Ur7fn4gun48YQX
PsQC1UYg42wHjafBwtpLgnBYLg7GaclP8Zep4NGfBSTxA9rF+M5BzKsf/n8WX9FXrdAwbpo8XKQl
1YkTzKYL4lIGcEewGDw6ixMdgWM511MH0OkUIoI6qN8YorAIyoduW17e8+dvaK2HHX09i0XNJaRV
beQkEWa6Lt9NL6poSfVDiLy+2ydhA5RoyuKilS+cHU2sl4CYFlZkU4Z29VidSvSKlZ8fzS0+bZLT
TGSvoTqrAu/zi0SzKy/j4rGSIBuHDwHGxUOnR30uG78I4UC/uYkwEB/Pzk9abEjBM/uaEr42sWJd
BCcDPHQraxjs0K+S20cPtxB/GuT2DF1PPts3bhxHRz98lNn+U+6O2k/NCE91o4iHaOuZu0v60PiM
wd3RDZPbC9OT/DIR6vBeORksNIMJ9Bp575WMdlOFnksOq41lmytFfUW38bbFvPmklQZuYiG3Fu6z
NPRfl6OAmuqAYqoJ6GdpUrIh5zRRB7sv1PzYxWO1kElHb58OyN8ERGn6rMEd/IL4Jmp/zcNhXimv
ET3xut5DtwUU/kDEM9VAcX9hZX/XLmYPKpEJW7lqkoh1sxLbDHq2NTgjca9UFgfJHr/DOytemEDp
mzspWHZfMCwFjBrRU/0gE/e6giMnlI+J+XiNMORmdAV41zvnGcNeYnIWFtv4sKqGV/AfRUim10Aa
lVnU5Shi3i/0yzs8q9iCCnW3l8bjgZbDkR4Vn/UpKA5C/D8+5WNNk/YRDmaFi2biRQm/UVPG+qIY
Q5rsfiydJLDHD69hqF3vxaAeBjq3tecNJr2mG4xlHcw5rJk1oxGlRwhyVH7pdfG8YJ+sksAEj/Yn
pvA0Sz8lEgpSWLLbVSqQMvJzGsJbcOvFJJWtgbMpAu1Q43UzffDRZXcvaR/b8o5RI3yjAF2oQZMt
47fSJKX93bfSZSfBe/pXchkZDfnxK62OojYac0HK+RqOKCYe2H0FSpqiV57atnmOxW+Iq7LANAN5
quOXP1iHLXIsSPI9jEHIIiqr5cDQFK8grdVq9UaS2aILet2nAwDUkGoSUdW2dfOwAd3+4WV52rrA
Shr7W3kAIxHmFTMysJ7uwla48as4npQDrfs5XOTX0lwHnWuutPRP/sf15Bl8m+O6l4RCJeZ3LYMw
pZTvKK7XcG84TYbswGpUhmR7x5Rj1BABq4Pv5AISVDmDMyAGqMKB+Au6RzvzFGCpsqQix6gTckrK
UdwjuXNKjIqezJB+qU/ywkp81uATTXUQibCRXKmD1zqZ+Y5fbpvPbtgQmzJLBac3/umgqeEMgSLu
0qq9lBBJMBi/yhBEvJkBtbgI8x5MScoe/AvRmuRvbqF1e1xN05jVs+jzRLbZAN0WI7iBfo5kR5xV
+drRf5/yxLK81Wp3udL2OHnG6ZWciqqAEEwSvU1bjHOlj2rMLpj+A+FLV68XsMKlXt0Uu4AvTS91
9jvJ1Dicb/sWwcfwPQEpg0J1o0AMbI3d6BxvuXC/nM7mq5YrvR0XifgoP5bbiQxrzmbYAJRu4zEL
rDzb9LXE0rKeoHTyvLahH+TIk6Ycix16B6SppIuwjbQFzuFcaENrfY/gljomj4iaJWkBey2WDcCj
wYN9PyF28QLBPYbaHFPoSRimPCOnwgh9u7+AVyKbS8clIDD6VpK5VA4S6asFLjdSXN2+MtWKr/V0
26dFdNI/WXOUj4StY1kXdjzdYXPpQxQvfb4VrZb7EH6EsnNfHt5CTlUx/lFGLwOhUQB4SQCFdMdw
VraUBzywE0Prl+Kd0LYhGMBpmCD3vWZGnmc/o4ixKTwkcK8A2scqVO3jkVasmhllgelhQIVC/4uH
QIYFee95l9jQoc97MUSUnxAEvMlOeQXznDxoDx5d8Jv/A1gd5AqeakaBjpFD1CPWjZpkx9kfaCX4
TOWYNPdT6SXvMdqUlCYckSPAveCwWV/NuzeMnCLUB9HaJNoq2O0Faxrw7S/HILnwEQ3MJ5owjzJh
FEsXkZNSL4Ay/p5TOAa8dJp5j9IMmoOVHCSA7/5UwUeRrwLsNHs4nULMCg6Cj7LPOd7NUb5qEQUi
BgJMntoWarsT4cmJ3XfUu16oyHvUel8H1ybpzysIDuZxGuoHHQDf/yfN9cIwDbjOO3EIW47Xhh7i
k9nCJhEp9RMaI82A5k6Zus0Acq1zqrtV6mhV/GGXi67WDwLvEffxW++WDwgI80RshCjSmaALsEw1
zCfA5W5cOZ7F9MEj3PFS6ZTxj953F6niV2P3FbI+9VBuztO4TEskW91DbC6WdCGIR34Advnib+zG
5RcsuZiy/YqeS37sZ96+H5iskd5Ih58Yzoe4Qlua8yUivjKMs59o/Q36MHamJ52iJ81m4YG/4LKv
qdUNQEQXgvvZyuPKesovxH3vY9fl2m5yV6oSsBoa2zJHrJm1oYvqDPh8EFynN37YQfHyStEyK5iR
bqcnzTWwQB8EYNn2RVrmEe/jPrmjhbyHGLctJnmMEijucDj86ULSyzJAb80hYFSXpE0Rxxjp839+
V9BDqJIlJ/dnuFTbTg36tjTy+RYS71+E/nVR0o8HwRvZbBSmoL0hqnVmLwzQgRU8KafgexN8ZQd0
8NQLSLRVhQlcB4KCg+LE2U954rGzHISOG4ZBHIyT+S01kVHUOlruzYHJ+cvjl27ohiamh3At6cxO
QbJxv00poxw802a7G/GPQuyHOYRwIaJ17kFEnot20BjfIUtWjqhWFZdfkW6mC/ohq25Aj88TgOAg
/egRjMBLW9/PFJTuKvnwSO4He0CHNI6oEo3AhJ2vc6sJhOTrJPR3PI1sVb61hz8NyPa1IpkEuy7V
pgeiOGxM5118w47GbdbBPlQaGBoXkNsyUWXz62yb1+158Gs6YWfGyFaM29v1IeRVN3yRT1gzNy4G
NZjg7WWby2E0TdSbaHcF8FuTBstX5M69/U0Acs1m3PI/hkqkpZcCUXYnq6mJEX/8Z9jfekbeU27Y
jJ/3VqoV9/NKD1kU3pZ6qWbq2euSz83v3K/c6znPYzv4L+rGkiY3Uxl/2NHHGaPYrH7sZM2IC1LX
ekFepuzZy3aEjKQ37SDrFJ/kBSP1ZJ/8+bxUTrlOxuL122WlfxsYMyjG0KyxWN2b0bDO2kXVfHzX
jONPx+Jp8974C7kMNRtbvyvARuxvkfiSBnY2Qkmi8DfuZT7S2EL9hheYdzq1B9MVTtzB7liRJL7r
vrWgo89R37h5yYfoqv48VewHvIip13/rQtG6sSY3SdX5bIXw8KCXmR5C4gCs1sa8TB/jqMF4bbtR
Bab1iOo48XIkN1yxZKdr7GfMcwv+fr4SMSA/peqPOI+Sb7LTdmGLZY2cE5cNn9xlYJYwepV4bfkn
GXyJeIMoNyujAgekDuxGuWyA6RCsyE8YKjIc9I3KX2YsznNzolGlpNIvABwc4/NnV2f2CIq51wtb
1F7vgxZf+ekYECnEAQkERM5vUC4Ch47iF5qJF/+RMJj45pYn8/byFjSWgzWYS2sKbLDnuZHunYnC
Jx1//Glnrlf8ONDJtA4dhryxr8gfw6ZM2+/0Xymqz/5Tgg4pBiYRRJLekFIMYh4TWgkQVqlv/+08
SXmbIuCvVHWjHvDDH33oLu+XLmVegt37fmKBXCDYTGT2gv1xao5HybdTNlLMjnR1KamBIU5UB1yM
LLCLDtWoDRspR96hoMemVlgQv+YyqUZwKpO3XjbTvcWTFHUAcixOmtBkPPwyy8H97DhT19nzDvF6
wWnjq9Ff/gQUIaxciBNWwVrOnbw3kn6LABllIAhEk7oVqAIedAhZyYONAHqoYyzQDxth57arr6Wj
H97dW85kPJXKOZzZKnXyRQGI2Jo7TLLh86g1PbQ2q48gl8b8KEV1PlTAjU50q/ulHzVHDY2bPxHj
q4Ejb1hdyFbZIF6poBWlS202AkKCs+QnGe29HyFGdicY9jJ6B8dmTY04ZYaiK/4SRFTUkGVf/0Et
bIxa5mODXbgdsja5lR8m5k3Hp1jFslYCp2HIaG2WDZQI2Tg2KvVDiHdIQL7fZMkGj7QKj4aRNBWU
Yuwab699xCjkXaAHUyGcuqIrd0SaBEdaBvF5JXWiOMz5J5qozWf4lBMmiXyGz/AQ/09U/+svqHy1
rRWM3M3AR8i76Q6VabKV2Zr33t3twIP25wk2ljNG/HfmfwRt7HqXF8h7Fc0NPyt5fvu0pwwajjJV
BFSkn+5jUOiTDzHJQvIscwiK0Medjasg43Eaek0N4xeHpzsMbdSLrdqQ3qNH9t1ZjHW0SX5zmWKt
b0qRFuxtQCleYP+HaIcHx4dtMzCV4dvtS/Ph5z0TfZdVx68OtP6DVO1dHDZuzr9jNBvensiTXlGs
MtmWhB+FXUlo4F0Uymt1lRsx0SbOM8eUbjbT4u1ruQVHDtUbYhGbzfdngcAfOUdHSLhXoaaSW+kF
Y2mETcTdKba0EQQAeWXD3icLcKCbW+wJCSH+dlkupiD7aYvPcm3ZJNZraB57RznfqLaETQvWtTbY
e9ZtJPeGJCIDQfmEjLjANM19MiGLn38ZMZ4BCJmsE/1m70AzpIeaq6ni9FjogyzeyEWQqyoSyf2x
3gko8bt11O5HjCQtoVeIdR6OAxJaYTn2ocdpu9d2Jhrr5wGjMWMdB2GAHcqoWVCHD0t/w8dTFTAn
KP3FHSJEAUnf8uHkPNg4mM+Jgts8m3llmWBcEsmIOKPAB9BYdU6xVO7DKPV34HPtFn/LlkUVefSB
2Vs+osb4EB4A0CKoXF8afAkgPTATLDyPgxvxjq7vRlnfXYAdaVzBONPV1cGN/x7YnWKbVq+s9YAj
mQ7AwTDqjgZTb1O7P+RadywRPp1KiRcCu55hMpO53rKeJ6CFB3IFLcQJHFaVHRHofek1UnXHJ9OA
3cj3wAT0xIN8yHnqLl0xUHhL1LtEzuExZDRvNvT0eOtd6o9ggbaboICVml4x3ObCGNo6J2R1TpRk
9P47ZQfgPS1z+SHPH+dKOPy3+kukdnhYeaihE82H1Xz3H/ZXrRMuYPqtioPw7z9dDWLQNf5pzoZC
CGn1mvSO4ohXOaQkGdgTtUn7ypZm5qT60biyWhxg+0s6inbCWDn0CtgpOhfi0o7YK5YOUstJHmHj
JplM6BkEXLlKi6HbYb26ohPYiF0q9/npXkuZV/cdnCJQboHVAihWK/+UJ0yOq1D8dFt8Q5gmzH59
RYmhAplQ9solPljrE7aUij/YyCA65hLGocXxHUxYeS9ZGtOCHyJh+ATjs1bBgGEb1VUwLicxSLRn
jxErqKRmK7IgOGfz0RuC4HwdRiSbdazDEH8hVd9Y4HyopoLgx33IVY6PSWwgykqAP9IQ4hOqQdq2
67AE90Y4ftC7sIKerJA1t/er/+JTry0rpLssU2+WE+YOfeOVdUR6CjmfKWp3HNyBiUZFqPIv11Gj
Y9tWRlSQ307/xEDBHXPlKVQePjyEgS0AbIfGE/zuwqVcMDyN4d3b0mcqZd7uA/p0ySEMsXL7Hddi
pCFMkOj/ylbOSzD2HLmE3492+xTN5UvHv3oofy7DPY1yTg2x3xXAaKYyrfOaH5tdYO1zAbCo1YTU
pF78vAfi/gZfERZ/3RCrGvV8WzX5GCV+bahKs0qmpeBXrzANJ9kVnEmvBL1XdzFdMJQqKm+jns1S
MIVnzAO9DfG6XRpZV2iaa/5lNFBsEePOL46UZ8epJnZAWmCp8yjH7UJT+K5yyBcP/lNaM5MBALdZ
pM6sD/lso7/3Ad7MEA1gOtT9HNU49Cc01C64YN0jN0PV+Z00DmTIXajfgI7ubC+qqFGxUcwEERyw
6AqprZp5AGn4vKxp5wMNdRMi+7prBBtjYb0tGvsCkKXHA7r2qr6HHfMVP4x3mjl+JLSS6ng8GXKY
EseNfyQRsLqjywo992IRO+8OR0iDq9sRHxpNgXpstaK5tx+kXU6gZPp6IL76E6L12vNVKoTKcMVd
bW6xZN9R34WKuk9db8Ax4xM5F9B24Ox1sXlqBARTU9d5O3bo903uMIuu1ibhEQo250Vab+xFS9y5
7Q4yjfM+Ucr0GJWvWCOmB8zjN2zAinCfPk4TRAMN9IT+/QqqFV2Z5PGrhiPAVweuWNIVH2l8Zhbi
jThRmhgYH1ABXI6tAQ4j/+CW8lVkfRGwKyJfRty7sCycdxfx1ggHvinl/1puqj4SOxCPMuA5xuK/
UVt8dZmmSQ6N2qr+INfrA4H8MQuHzdaraKjZ9gSYapBGezRzLsWFDPcNwczUUW/f3N2N6eYlNnSW
Ioq7+L06dsuTarQ+YYoY/aA2bC8PRGpt1gcxJCYuwCdSUeg5pJFzXw4c0oWqvqn8dqizR2ZIg+oF
IHlElJxGshozZ9akgOINvFsOW3UF496pQudIC/mtPZKF4KOQ6zvB5XdBLOtsQcLFj1TL5FhHNtHr
+iSKKjPkh83el7NWa0YNOhlz0QtG/pHZHdXIJ7W4nmd2dQ8v8QgpPLM26f7wwR3k5+vXAt/J8SvL
fCZfzb1oGVZOLbTlWn9A7aCvPSf5qMCyc6F2fEvRoSiYlMFirLGo09jhzVjnC1jmzHMOFft4vwAc
LsmbHfqVrBZ1mAZ2QPDg6l0yBu2pHFuKZECMbxm5wMo0FcL4gpKhIfrADbx+an513qFlIlqbGSFu
dqKb4ItMRY8AM65KSfN8FAKI0oDd61jBHI9ijAReXIBjMcErpv/vY/feT2gBTTfdvnStmo585243
NYrU2as36qOdK4LYaCHIxQWJDtNt/V+8FZO3GSY34dMaq8DWiwxB3q2YnFrJP6QVhSOOBdai29Au
9nXGqmRsIp3v9WTxpmZYRQHK/oFaQfOHmBJxv93RBZ7R50FmOvlElVOEAWXCNN3ZdqAg0BRZG83s
+uNv/6ApsIMhF2QuI/2XMud73E2Y3XO2hjdR2HarSfwI4b+281Q15IqN28Uyc2ckpV7c/UhG9DSZ
+3xyud4MwEpKiE5bR7MO8Q+AY7dxEcVTw2E/uvnkhzIlFos4pCYE7kGlmyYa/Vb0VHiwDHpyEuOw
LjpFLjnIzpphm4LuyADjOOVK/AXR5zo2nskbaST9G0A+6RoWLn88XtUa7+YNya3mMmANUrZSlslt
R848lNl8zDeQYVvolxt+UYjRAbUZ19xyjU00It7S4C/vOiq1tRyVFW6B2acKZyQ6oGZ+frL3/CEW
D64n/UFU07nnmJdEjf9oOdnyYldJCztNSYx42faSluBBKit2Dt4lg/UXQ9VXujR6u6NtsgcwKTdI
z0ZlVlMbxLLCF1LbcTGYjRYlsWCDwjBnRoBBPeeSov+RjGuPdMzmzVaHJK1DoR7drnywWkSe2JUM
X6QxfLjdXMKwy5c1CmEkaRrgNabZnzEii8B7qqXGaU1zFq1kn/easdGeq2eo0dBvFed9I3NwUx7C
fghcdxAwjmS4XM5cRIzXBwZrPe7drqw4xL44aaiGfZaq3eEKsqQq40oQ2jcIqzU5xeKzzA3toTS0
xFzufMqy4rRN9nyPqqrFuseI7fFPCzA/0ee8P35bhlN9HfmNEA8gGDVr8XaSo2F2eZQKX6l3n29I
dr2+ohwvf5jDXAkGCScCaxDfqcOejwhCrOsV0FTrMCvW3f8yH8U87z5GS9bs5mta7MLXOpFncpLf
Q4Dwae8GXWZIyxZZ9qMAa7Ndak4QnPbtUXbn8DLFLsDA2dfST1z/saQn1j+QWVe4kytBhAOkbcaM
bEoGlPMJ2gDmg/smb27yZqN1sqYYRFh4McyTdzMRENZXzAcIIh8kAehN/S4AHUuINLetswY/BsXo
Mo2IJi8to+MeVln176iLRcmR4yvQ/KqwwGbpwrAHkHkyLWUwfjJOmU78gijJbrGFFa5pP6zkYNg5
FXifsDMvj6HFPbkR2ORFtFGt44Ctm+HlAibpZPsel6tr/OVYUffSQUO3oXNA/mYhiCSTiAqHvsQ1
BcE4P58GDtXRHX7ofLd7eMobHVb3Jff/sq8cRyi8KlJ4UcemWr2ZSN8g74r7RUDHN0vYFAWS8c1i
05BwNl7fwI5KaMySYMxhsYL2OMaIOBF0Uza35nqTzThpzCs3+VbiROyR4LJFHxiw+cHKZgeWeRkK
O1XUzThYJtvGoClz9B9q7gVO3/YApf7uXcg2XxbWeFEZ+6YR7OlTHUXOH6qNyvmYbbMTIWc43D4l
4Fn3m6xPASDIiJ286pPJxRBwIrxe9IuULMi1Ax4rVqsBkaGy/k1GPbZxftJPZZJjwhYuvy2qjF5S
SG11YN00WVtSd9d+0JM4vVt/9qlvPxKv42txX3BEWesYam1c62rBR2g2wHyqdf9dOGFHagE7VuzL
iwjS7ST/PDKOr2MPfUvqkYwzmRSil1AK3mPyw63MvPsBrlXJTACl3R2JHD7T+gGlxWuCx8v4+EKv
jWvDdSqXWXCVrTwwlrqgQMbV0rbPNmU5nj3nF8OIHtbVdI58FjqeA3F/XhkVP5rtdanQ43ddRwLw
3vuKYrRt6q2A0FtPoHKlkTB+/SrnIl5uuazpB86d0Zfh0q3IrTTR9YFhwQ9Y6Kd8dKyVX1u9Y41h
IR4Z8s/t2yql3y6HqJhQj6usghYry7vRTgyEYzeBHH1FowOYzw+hN7be1ThwP06Mc91z48gu5R0Q
QBfi8Rv/OuoUF2Wndh41IM0omncUG7rVB26FS2o1iAOyg1Sii57n5uj71Bl9IhXGclmq3b4epORs
fOSKwde1d8L9IBEWmeQ3rPfC9nH417BX8cXiHW4EpD2Ty9odeg6liQTgz91B+9higKcpazrNirn/
EUvXu/0UE2ei45Hhr1QtfudctNPShRiaCSXPPyQRrsHWChBz4hgkLhSSfAlSHPp5MTn0k6a+0zgP
y8W7/3/nMZhfoun6811erlCTmK7RktoxMAGQQZaGKkI8SkspKZew/BXew9zgDhvPRPKNY+d7wlLk
rZazxQJ7Eq1ab4kGljxnjPTHzVkc3dDZ1dx4vaekP6X4E+hcdmnjNv2tcBY1e1K8vAAK1LeawCPS
6jYnzZcHMPpV7tRLemQ605/uMEy0onRp3+EmP3dQ4V3TzTRu/C2d4RlUP9fVDUkEbkbibXghrXX4
ZWSRkoIEdnt2mf45f2lEQNnBsycn9xNGB5MZEWO5iUQZo8uWyyVZ98ReDR5eQBZqOnrYaelkSS8z
NK4kEw8P2e6/8LdfhiVZkBsemeeI2c+qdW//IAc0fkVIS62kDKGT7En5i8drkiZ8gV7ymC76TG5K
3uM1TMzpcmcnofs8u6UIEse0XupAn9RtGf2BANQEfD+/lY9hzcGSxcB4femfuz1gXTJ0k7IemO4M
EtrqoIY8Ds1iZp1CECTCmcilX+5dP3iNhR2TbKrdhF5pqCid3vZ4Sl3FWyXikUv8Dv7w6NQlOrMH
AIZZIAasDWVon4LoNC+6VeM1cSZ9DDn3oIdhd8jGVfUoZhU27w1lVzzPfTFHnIvbzwpWFk710CFb
7uYAZn98hF2dtx9iWccSEsvoSUC7xeZ78h18o0YSivYjGBcjEM50bKL9MoEgSST8Ftpt3qoLv0JR
f45V7gK0Yq9ewo/7/X2IHVsqBijJ8oVbeJvGV0xOCJLoZyMSTDepyvVdtvtB2ORHST5kWOjTBTAl
w0aXiyhDK5+vsmlzGJsJ8Z1ORVIY/44HXSBg+Dkr6DKnZFojCUGZWlhtEfuGf2CmxqeHeuPlb6dF
sax+OFQGRxfCasUYcUdhfMw2aEnL6M3uZarufNtRVEu6KmYxi8xCjL9akBJu0FY/G9diPM36L1et
gpWAwUSvUKzr5AtoC96kFm6mydQ+G7Re9GFR9fTHqKQRpbiMBpAqGSNkS4Tb3HDhShsuNuCTZyUi
Dds1V5VsUvR7kvUB1sV7l+6OGqSVRKZbHheyR5I+P2b+6Yka6mlzwOb860g87vmIdyHeLoTNSK6J
Z+6GMq2sunW6eHv7ZOwkFrTzYrACooU1/N6GVzuhc8xtE2NltNeLid5papSdMLVWmjvhBGjK2Oe1
RUg6GFL5ENK4vPbfvr2Ks7AO0+BS6ZmEnB24TaQ9TgnFxSOGKpWRnNDwFRHNFJrcEmkpyVZYgGD6
7lKOBoHdAsgXGPAC3sA6bBPvMkgcUGpXIyfwa29XeV5rCzxrsZsnh2mcqPStnHTNU+NxlL1qw4dc
vK72G2424ghzM5shxDP2f9hHQLGceWaZPiSBdNFfbYfWzqyhvJUITzdkDkHL0SPhjzPaRfS90ASr
nuCmwBT1Jz11aYrTvHEGdkR2Zz1EAmiDr6LUWK/ROEoTO0ZiRq7wtGKntTGchIgIG1loUJqpgEXO
bFW7rZUIS6+jMDhud7+md+9AUWCpXS+MmYgMKmcG3y13SUyjT5j4sT18p7qZG+MZjPZ5Ew6L3R7q
YiF4kbAgy4Q9XG5O1HvPbERh/ZZrg9M/prPjMigTSiw+W8c20kS+0VAEaZxoc2TfqeVnH1E+82Wp
hpITv2cIhbJbUxf6yRCDrv5JbLjPnfENDlUtDibbN8zXFu1+3SFAMpmyXN6N36ECpTRlvzg/pFP/
F7KTap7RwVl26wrXbUW5sFMBgddHggspIXzbpQSDORw5Vd/9g9N0Pb1vtPXGThmVOo06XBJv1wku
QTFSLrODj3s29Un6C+O6zh1/aW9pS9tQfTkKogKcFBUL0JAhmqWEQ24jjNBVUcuuDsI0i4CR0F+w
2kpjRZRbhcqwKNu2OW6KPB5+lPeAHzdLv1DlcpqVBOltZAjIGzwkPqceQa4pr+Z1Uts53WnP25HB
h2FBQXizYHwEKOtfGLhi7Hh+eQ73bn1nsIbMQ+EMxRK9++Py+irn8snzbUE7tDTzeVUZfuZG4Z3I
Pc5xBRVvsVhx9WFLytfL+OreBRZiQCwgTdjb9M2t3YtifRhKVOk1e+FhkHhooZ/vUVbft/gIvjZ1
aFTOQU+DahGcN8jusyzc2xcUN1TI0ptDHHshK71Jwvi3y4PQcHlS2vp3eqtKQI5UcJGjldQg1ERm
wnv+ucAzAAvKFNfbat+cJPAAhF8Bh++vVV8YLffNM7Y28Lztajjjdsl05awZjL+v9gOkMpYLB/IK
SoA8h4zZRe+Dgm7JLszKkOT4Uy/aF4eiCN4f00cdbyH9ogUiNhGaT2fRxeJ5dvCA3KWsLUk8Q0bG
fHT2u8EIVTmVUnTegFdfLTcmDm37VMQqDFB0paNjBhXrZDSMtXtQvVKGt5gW3AvaQk9L7jVr5V96
pojRXw61ijY9aGKVrvLXVJ+5RDdIv0ez8Mtv1tQxjltloUZzDQsiZJzL340vx5ASFU+NPMHdypdn
oQJAer7LYoXhi70vYqUBsCFGFHpYDy5iC6EY1+H20JpCNqjPqaI9rx3KpUN1d9BsYiSXjjx2cwWf
dYbm3Vhgjki9vbSMPfP7czS000NFypSZyl9NRBmfArL3anFjtLHEaOFLIn47pFq9USTIY9CYK6wB
kv+RDDvLK2LVRiCQHpchLLUT5AsWK85mmo+XzlqBf4K2tOvR5WkpMCo9fcUFoqqXmSBHAWbUKCMg
4d5+dQS8ENxa3LZnZuuA2ms6cDCxSVJjng8qof6j4u8OW0T5yUxKH5P9TUGh0MeCumoVZUv7mKWJ
/FhPdKmRMHEFkkdVzyqGbtOdv/8pbRMAq1vrxMTGvrihxZgRu5tRj8XP+6WhaqfM0JDu1oLeVZp3
hilWAeZARHmJYe3idCa7Qpu5xapkewmLOOCQ9fwwFI7yMS3saLiCUbDDggDNh5DdQA4sGJ+KfIWM
HFuVUglLoKSYc76bPfdVeAEvWkqnM+49l4Lb6w086jlY7AO9Dvz4QItGeXXRX63aHWHtbAjXjKTw
4ThFLoX0eWBTrnzkRTVtMYv1xdLjm1LhOarLeB1mLaeQ8hB2jA/jPYO3f5/ZyABk8p89/cNNKtG7
te/K+2/oVa3Ev1bG+f+6nU9+Hl7KE4bcTi7bi/fYM+9v2ZNmGAL/fnSLxAL66rPj2dpBaNN6N/YN
gyy1h/8b8fihIkHdLtcoF8/xD2sX4uOaVhqqW7Cv1O7nX50Fg1xaEEEMwSWkjkQEDL/pRk+h2cFe
AmAVVioESQzoQ773zQAXJ7+7NnYe9ZAkR05FJWxPgl26KUQjL6mPOv9cRw6jTAWWmkz14PkIIvIQ
957VN7pN8069JR1BcV16OOEuAcfPDZk59guW1w6peHn1tuJOrc7ZTXXge3yqgmseh2HdGzSuj5kN
nokh8bZuFQ2NczkMO20kAs1GzbKaaJSsQFhOM26udc5iqaImi4Yo+RQdhD8WEm1w0jRsC6MlfbUI
BV+lVXAqfZkg9Tp9jf8P0ocgswjM9Y1mH1X5m3Ji3euFh2DQ5DAdWp+MuqyOTLkCwnctcCjEAiOm
hbJHGJwBWw5dA4UevoZdhNLJm4TggIp1y7o49wG/lmb4RsqvHEcfHfwTumWocnOR1ZgI/7wk3JGo
4viYhyd42/PGPgBJ6I+aIBo0pYhUm+h5jx9jmNsJyjssrNX6nyiG1KI/Zkoai9BYoglIv4vZ3+pK
Uhw9A9LRK3ZOuivaoYKKoBqtHYxx0/O+ZMYCuXCEvvglgR9bwaA4F1thAfTgmRSyuTbBGaevne2s
o2HAOxWVqTNxcvWaHib5ii6Pn329Ul212mCF6MBndXZGN8ORkw5XHlos+FtJpmHm7NYQBHUFAc28
5xBcp4P8MjRypZm6L06XYp6UjOJOXCwfWEryw6dh5CE0xKYlODQCUf2EuZGCfftlv7qfkYqmdOdw
6gkI2XIiziSa9+oGEs2FtXzO8qjcJo5ffYuybxl4Z0Vi0PCsE+vSzYa0t08u6pGnW2A7oJi5bLds
EM94GrBCLA2Jo1UrW2fUIO1MLO75x/rW5dulsmzNhrqIGTmshfIcg6iJ4YlGozW1ZbsJo5dt7LU3
DaDI1TGUpIoEOrwH1/9LXcP/aGayDjxCMLVNSprvDXqDrmXD0KAosMCWVTcTEe0hK9twvRmvbMaX
BhQukyzhGFgyy76k5AoVPo8IRkvPKBYoXaxAKb7D+0kxwok2uRVYh9lFoKNb+CvwS2dXidbv6KQ2
NVLxYrKVKWGtxiJNpPRD1jPEGBoZu9vZPxcew8V0/LwS2py5db+T+eUVZxA4/932W/C8x8+PuoIr
2mMtY1yRaj2yL3X1HS+Z5/r00yQZXB5g+w6bq1SE7iDejAwup5hp6guQfzXtrw6CFWVSppo2rDyA
eXD599BkqQR0geB6oXaKmKRAnI0cVdNjwesQ4loRst2GTzPA2hFb0GBXlK/22Q2WHhKUAKCj+zYF
M5mQPY4wZOsBMQFOk98wu6sg9NE9s7UpSsxEjEfZZyf3usJDzo886yY5LPA2TqGRe39zDJNrgNvW
uFPdNglcu4RK9Lq+Kwwu++QgBDTIzmAfVFDyqqKy56eTxpLS6RqE02CPYLNcFEAxaD47XveCnZp9
iZMYjrH+2Thv6aI2IsV6SOhiTixWPaJrLDKM94Pp7ogA46Wjv/GXwXTLwHE6QuviU39aPcPDkUSg
G8BPc5xesmqZZeBb8it89hjc4ZngCGb4KoQn6kv06o9y+7CF1RwexDZu/d7GJm+/zJqWfnqxnQr6
HBf3MZmCov5Fve3gCc/toravb57UIpVl0nku4cDUNP3dxWg0v88bO1LYDcoJ+p5jMcXlF8wY8m3a
y86LiJD4N7kFZJtlEK8JfrHul3RS2EGyb6vkkiIFx1bO/8oeEW9LTjdTWB1mXp3wiGhRt/pkxwGR
koJCFh+gwu2X/VcCIgRkoxlLn0ukbvN1iljZj42BAPwZlH6goPjQZnmJSy6pLw4ABaxIW9Loqiih
pDHv0JYliTrstkWd5hVgESQ3ovudxnyotOket62lqouhIDZ0WBKJ0M6ur0tQIBquxnmxirYDMoKD
rDHali6pcSIjGM0CJkW5aDUBdmhYqSjF+X6mZXR1m1KAfmgqC4OD3RaF4QevR1uWieRGnDMwEcAy
5Jh/WkD50kZDQt51SFGwzmKmHu42igxRAwG8U3hfrtjJ3TRFmV3hBJT/V3LYcILeGSIyxl8t/1V3
//iGC6eXW2/Poq+v5XumYzaXI+plN2ZBejQd/clMVjiTIAjoF4ssW683547Pf+6wwZ0bNlfpub/G
vqCvLDGtrQRf4TpDkWHCQ6rZ0H9XLtHmcyYJN2lMF5okmYbdm2OvF5DQOo3fBYnuydKcFIkFYEYH
BzQ3HG3p8au0P4LecpOP2JQFuVWhVdapmTo8F6HfOZBlTt8WwaG629e0YL9oaC4ZlQCVhhAiPRYn
SSvF3Y0mJIwl415aE2bZLWjo49OA1WA0ceUXMvTpY0frHcN8yoVEGO1dTd+86MFdV8Scs7PIX7Gl
cYue/FyQDGdAA+jyA9oiLMSVkSBokZdaqJoUybS9TFkpSmyomiotN7it0GPaLWoHY0gu4vHpr1Bx
zOICGEKYtzXjeV8OLyWKAFOi0nYdKcU93CzvMFlsorhgrd8PaTXv7pzcZL/r/OmThGMoEF4NOD1P
JkC7X7ajcPAb/VN/oAp4Co54jpl7QBe48NtOn/D8sTHgSJPVMPbStuRt3p/kc841Eq3jLhANgAbR
c212CzpIW4b3MhY8QQ2f5AIwP5tx8H+Fj3XtBM/iojkRQ7BbbJZJyGSE5MumgJQMj5nB/Ccs9DVt
PI2QQUeeM/T7pKZtjEndyV1KeKzlJag3JZQvkN1yexfV0qJ1dnEUptFvwsbJB2WHb17fTii+DNJ8
NH/Rt8BQn5FsAth+0YoG0RXZCmqrozKcXnCOG2q4jPp5OHy6LIlG3Tn8Zzoi3EdRGYf0Flljh6ut
Q35fTAlLxzWUdPsDcelsSikv6BsYOisw42kL7A2q9JCbgVqTPxKupEDa4AN2l/aZp3NRaCWngXLn
QoQ2q1vXmjuqtxYFjoz7sjxUXjEidt0dZ/Uw1WeHMHRj9PoJi01ScwibPRxE4wMGgVI7XwmfEfxA
SY2IXUBuhSVmzkq9sGLhqZwglW5bCX93PD+V7m7NRVgUy++awFHf4lnyp3iQnQ+MVxraVoVcFhPs
MXtWSrWnNsiZjhVlGf7e2WMW4SKOiJcC9REgEvJTNhy3Zg1UZawJeB4Mn39dKwN5uW2KGYteqehm
FIN5w45FLmEw6VCw+7K2Nn1rA5pAostZP03hy73GwG4YI7S0URksFapdhQVhOhCTC98k3oTEhzcm
Ma9WgEOnQFEfKzetWth1TR3o28rlmJG+m9PQgswEN/rBCY1nm7L+Z4gTXMoKqfQvbh62/1rMc5pT
AnJ1TDiGFejz4cD/4srhoOSSCE1JA4Fp9JfxEdWOGh8FdMys3LCUGn3ZZloWLgmuwijTpUSO/kjg
WCs9WgIrF3TDtE/ykwLMDlEqujmfTsoBDdqevYceALlYcTWj0iP3OdQVpb2L3WzNHno5ucSPEjX7
z2N4L3ndeispDLqs7SI422LTLIt9+X9l0AHDySL2rUnxwyiICVAUTuxin/2j2fnaDoI/F43i6HlY
S/650Fu6sgmSSkDwqEcb5VFLyMQ0NtxFEqwK95vl4zLc6yFvOPs7TEEjavixFeoWddaO4Rv/IjoO
X72/RoGCI5MPXyfXZyrQcExYBS5ZiKHzSMueOLnh6LgurzWJarxVqjaP5q1b+NH6KRoE3r7tcf5I
JvpaKzQ/3Td+yo/bpOlIT1Dlmfw7bJronB/5jnaaPKLs3q98ZshPA4vLcvAuYr2UnDW/hBRHomPo
QDi/YHVdV/D8/pyxLHPUvBaFoh4AWoDsLHKzxdfhsLK+GsJGliMsreoCwIOYf6u4yY8pqDzJsrCA
rEeik93i/FUMqolqFOr5fxjKiieZLsQnqUL89YMuRt8DgXtO6IcH/20em03u79kzTNhSP5tzOqQA
TcfShT6JVVXCMuForCzO5DoVbUbgHZpkfYvLRKqZS7Xzi5QLxK4la+G5L3+eaWpDEwseu2UGn4p9
K79fYcWk6oSFgwlE8aQpwrG5j+smDdUid1JeEjcmAlE5bfBnkGAUQ32hJO3DN+NsGskjD8Y+/Jdj
pb3/nDMXa5WMbqk7RrXfaij82VsVjwqjwzhO7j8wih/3IIaOkb1iihBZ1/Iv0EOmg1pjRI7YMEPT
oXAtPL+9Ws2X5z3oX/TJSJtpbksP2LA1fkr/H5Daudjz1vDS3cxCZGt57j/iISV50J3fCxzTJCnw
27QNsJ7eww5n3LBAE6GvYTeEBjKrAjN18RIEt7LLIZovxali8foApTECXn4tJMgZD2pP2Oguzdsz
boiVohS8BJDl9nIO9HjIEmsUnmyUFyMUZOBnfuAQlcXhdkXWDR67UmJ5LIJPPO3P6VSlFJRFnlmr
G8XfAZ7M4o5rtOEsxOqlpyyA/p4wPTCZwUl7O1gNQrCAxXHv7guuoMwBuOItiH9bHoba+7ogwmGO
Xmkq6qwB3U8YuZg6Qi9Lnepf0rkhdyHDQJJV1E1XYJZ4DMti18OqgelX5LcgTF3E6m/J7MwiWTBQ
rjFaRYMPQnUNrjOG510q9Uo7IZ44ypeNkdWR7jYmKuU+hF6O2TnQP09LEJ/Ri02sLhl2gVSDAirC
v1x/1TcGSOXuCDh2QiZc75PWEI/XRQgeHX+H8ci5SmBth7LcpuMyR0wTdB8KcuLGGZpa0UvwSh5T
oXaGyMw8qZaeF3U2ABHkE8iONRx5bV77LjYajjLNV/aXsj7x3Mtq3EsRdYgEYsl8CITMIDxzA1Ye
TPsPZFQRDQBYzprkRgi0Jb/WSahLbzbeYqvGMFyoWkn4wqQeCBRV2DoXjz28wsuy7zi8kqfEE+4v
ZSBYRHeE489wCsFpD5syDNloCulc5CnHD4baK4FKepRS1dlxHWED3ptd1D5Y9wX3akSh9meb4Mkd
cUtvRBQVYVtXbx5hu80Bm1ttxdfVs/mpes2KV7erZmTnGeI7QbW6YXCR5BgLpUPZb5d8rlQrBmf3
rgQmfOaLdpIIVxCYAR/4z5vkX1AXdX1RDZaBbCSeHWI0S0HFvpmM/AJQbRo+MONyazn0MU3MVkTP
ckVVoOdbnqxWLlzHqiNTYFZCweTxFZkDCkQZq/PFkx2DOHkCn26x88wcrVpxLNePMBB35BNNbSZ2
7JC7SKSShNFjOxXTHfd3ZnAm9XODkT8lXnAVNgJo1JZ6Zzh/azU3whUMXwhSi5pWcu67ZfhzwmbU
vK82UoAej/lVk9GhOWwDjaGuHGfIrdKKLk/b8K/voTeutK0N+txF9aiDp6PldqNHaqPJhSq9AFpF
3NlZgCD7Xl2uckZ/lhmz8ZvrvdJNuxwU3knDGWfmyjE7Sf3ewfiLcTIBhIGtWX/kWVsXwekpNjM+
XobHbg6s/LcZmF2A/wWtFQJGqYTabBkPL8rAMad8IRqlVb+5o9HLPFscm3noxZnlUGqkdNmaLs4C
ccZ94XI0RNgIpxNrF4Qp8k6tlaTBUwmbDCpXQiHCf1ZNAEakaHzNUvhGUvw74aAq/mSdih45lS2Q
uU12fRzAiUSsP6J+WGXK8NbUA9uWGz+IaOj4IMHqlfb9i16jOT5S7nU7Aq5W7wAcUyjbOcAmochM
IZcD7+pn1pIG1CBnzG8sf/qTU8XV4e1afwdCPzeMTzD+QS6ob00dsEVyomtLprBhVRh+58mwyq2R
MJge9Vgw/efDnDn00m5FEGBpk3DaNxEQCUv4cT+wgZGgTR3ATYXdLLegz3wotGi2XwxrZjGPrW7l
G5zYvXlRkwtbpQN6w68O/IeHZ5R3ZGqJvfm+xgzqpV9qOi4paPsQivu0fC3+KPHE3ebS5Vjpdawv
1QOJ3z3hDltqKf1Ko6K/7h89DaA6u52YSxQftK9tvMcKvVZlZkqHzwe0ER6OGt3WUuoxENswN1sC
qQ6NhwHAbyWnYcjE1jlFkp/Ape2MwTU0hQs+nU3qaVUlqqpl1gK8/OKSu5zvNW7eTvAJ34JGTOHz
4qGbinqq0nEV5qFLBO1PQEdvycgSBPua81SrrhAP8UmJiNUmpH92T8sSMXZY0m2bv9uhnf5yow+X
TXjMcya7XLMu1ijAAV/DgjHfnuWXviBjRQMRfnFRCuMJW7s/ZrnL03zciLZmidXgo/YET6IP1GKm
oWG0w4cq6GWaznkirv8hc7BM3iw1ITVsFlJ7UK57B59jq6OjGVhcl1RjQ+I/Mdcbq4nXU2dfRaff
46OddI0BCpa0MLmylCx1CkTan4Q6HJ2CJcoXuY2VPRHcZo+UvhtQC4xZ/tK/BXOkTE2HtPhirR5t
QTgC+7p0nGBS/MKCdf3AgNKa20NwUEctYX0IyAmG97nAheWxiHYLgpJ5iWZV6tjq84PYPOTUHb4R
Dz14UfiyZ2DfhsXZj8IEYg2Z7nxQvnoNXeA7XEandpCW6VfvOtXuBBr35WKeFtvkLMoAp5n3mRIR
dKQbPhkPc38JgDsz/RhA862ymvuoLbWhUxocS/z1v2Y6ZmAOYDDErYqtecPLI2OHF+XAyX4SGs11
QkIhz+HFzS0tTAE9H+aSMuIkeHstdr0NQexOPQlqrB7cXr/lBs8xhQckstk8Kk2wTNTtjmqUyBUP
gFvGqKCmwLmMNp7DYM5cTY0CgsxT8KV6KDDcObqYGxyTyUSJEcQlWgVfYoJ5TlxWFr8LQVPIJ0qg
CIVHor7O9CLtXYSs9hAmz/KxpDa6AxCiIryyoZKV9QYi8+YGFhTsr4nAq79HKhO8UjHoeXW4UzbT
B4LBjd7M62UaN5fWmNNNrNXE3OOWkfUCzZdFFLCADNj0EBEhv83Jc+bc1w8ccZv3qX2MfQfI8vFL
xCHDs8POix57MqBuQksvoqZ1RRvWyCj1j2LdN75tOul9IIZOByTHYeheUy4dqVtXVO1Sa5bjzc2A
7JkZ1V5T+hShFnlHrFa/nGxsyajNnJB4j3xmFTuZ2Ol0/wt6Jcv+QqlvKF2wzutuqEHYLKRsMY/w
2Nvl/VU+cPb9gzuJyWdUrPcMxJ5fk/JzPefkAo2/2WNw/5WoIwz9e0e+bWs9EaoauwCLLytaEJ3B
lnsk93a6VOGr7NSR4ZVEY7v9ZQ81BEDUSB9kn+yu1RC+OgG1s4uJvS9L3cYe/r/mFewbQV2OelJm
9I54vF5QiaeJPB17Fehf6fqUPSYan3vidsch4Qx2CEhONif8gmN2azXg5apboRhNnWggwKXox82L
gMH5z9bU+LW6kCyxh81iWl8se0RwU/+i4ZqBvDXfin8MFnpdccdgC+g/yHc7HxtupYw3UKNznwSo
DjU4EY/zsARdRTlqy7ABxnCUeTpxTEbVlg7rXc7/8Fgt4NNdGzjjILh4ADz25uKePevCtq8Ht5b+
ZccDzc0MBnl7EBIKLouRHRjKJIhizMHEeWOkyIm+GgezoY6sqJ9Zr/Ztss1Fk85RymZzmKOJmy66
CRMXtHPcnNTibLidXJNBdXI+65nN3GOKTLryEzqDYUZm/d5aVsyNzlNJIQB3/9hkHec7DEbwYPoK
fydUBRre1/PcyRyEAQFQFua7GA8EkPl2ChxrwFQa9L3nzPAs1agkG0FSIyLO0E5sqAbeVm9BWrqD
NLcJ6GxhsEP3hKIEszhw2HInc6GtzBU6dRy0vdSvRgJfjXwLfzQ0LKfL3H1W637KYF5ueNWIOLgb
LSowHkJpLcHW+gbWS13pTxFqgYn2IBxjNKyel5Gk+CKvh9Mzg3Q6hRNVpBzFElP5nIjQeSlWguds
3ZZVke5zmVRB9SQg84AJrTsBBV62lmgvmdAYa/YJc8/r5BulDxJ/mYDrWnwX/K0W5FBy4dueBSep
F2DQwUmyiBFCkSI6XfbFSX4cSWj3CXQOcIy3/8vM7zkfzKnnbyxJ9sOl1RD1ZpzGnPYSFrbDt62r
ckx3I/I3j5QA7IydJUL69RND/vFzDD1lapmwlTducfMzuRaNU4vlgm6Um+cgVj4Vs7spQyiuZLB9
seqeic3aD5YmCZFneq2yLhu6ZDYId5h/2EDuYpODlV66zxXnAW/aH0OVU7Q6zlxmIvioS6R0rf4Q
ENGdhvde3iwwIlk/3NW6a4IQllTjpb6HTg/n0aXG840jUrkGcYA0rCIIAg0p+fKpuul8Wn3KU1FT
3+RiNCIiFIPANwyCKazs5LkdJajFGxn/dyEsFJuiV0KgFEhmOJSWi5lik54nKYcnje7Yqo9YXz1f
doXX9A59Kk7MeruaviU+RNoxQxpIxj6eFvfmD1QGgKppIh/IGdm2AgQm8Ylob/MlIy4l8Z0Qbs5Z
Rmsqk7iDW5TAa2jILBFNFF9EwxsWi3jRTmmswmH1ZyDIC8HKOHoU6ONhDIwB7Ha6sIkibZ/DDquj
kRaXgqQo3H6XeeTTeMKl/4G1Rfyxj3Pou7BbBh/5HBZ+/MQPDMkvaIYXvpe1fN+rMNUY+jJ+3z5g
GRpl5uEyBZ5zf8ZovRkA9WegW6BagFwmDhapDg70mRILZU1bfqkNPt2EqWzH1Pdj/yn4QCPxAAWT
rhpHjhivqM85WNsPn553hpYD+cRrikM9aWD9jTKXIAwVSx+0be3vvH5XdXN73Z+WV5D+KB4SjYRT
orMEcbN3SThuJotLECGZ+WKHKYrth0cN5zJsd4sTexKrDoAgC76bTegyNyWrYWc7fIqc58dpH7vw
+tc7lbe1jL6oKj6Lu632OmrU+l4vspojPOopJor3il8Mbi7Fe/86Jgfv9gIHSCVN1NON2WxSm0Dd
u5xz5MWvO7BTvXI7RnNV/nCEe5qmQU+H3czypTt85gNTy8ZsPfkNlPk3wIXDp51f0hHC0bzJ20D0
JyeK1hjZeg2pSvCA+/rwnX0pOt+jkeIWF6xVFm0MOmB+knyQHB8AFpby3OBhlRP97OIacSyC5xIg
ohlxZZNhiPDzTrQS5eza22cFUyH464jyIcoxRRB4gQy/9TFCYi2wF/eQhGenXVD/NqeADdKG0Jej
muH0NhGINt7R7X3wNYG51g9HYeLcGlJZ9q/ESNPglWD2QeYbGL6fUX9so0ULPVhos8xd+SoKbPq8
LbrpSmaqXA4YCxEgAiaiEnX0R95DR97CeKeHTRQB0jBsT76MtOnNTRgMW/NxfEKwWGcCujDRHezU
GoXE+2grkt71jIVu8Ev3FpOVv2r1XlX8h0WKf78hZtyrJqFfkxDyXXHnG+IXxNYib3kjIQFP88Fs
TJ+MZqoKXLvCG0oLsjcCyL9Olq1bOMr1pQYYx1jzkHNItR1kcsKbgaMLkHNdMQ6UqSxXA1LMxiM3
N9prDs5YujuimM6C9Qt+C8Fb6OgN5WvxDyI4FJbq5MsTD+7qeuQbsccAgwpa/036oL8xl5DExA3o
+5mQS7qqBPQYwi0yrl+BkB5qUGm/9VlO3GHKr5EoR4hOty+lYiA+pQlNgM8wDInI7FNGisYUmbJH
FM6SGrWH1vWl7qiKPqwI6Qfj6HcqI+/RSOu7HXHrEdkhl/OrC/aPZ6DJ0XxJaeB6pb/vb4/Eldwd
k364czhryMum/ijY7ocSZkzBqiZxWX4krW1PUisnTqMfUPVE7v/dHd2R5MVprKB4m8CaK2WwXnhR
uCcEg1MaRbJ03cOru2rHs5KdzRQP12Id3/C22Qzq1xBcVOrzfjozIcIDaZmkQtgmLx59VLjsuHNf
b0BVMIlKiQwApkHBALvv6O3ao2x7PhHLECLTDjiFOmBcxqfqqOaAGvEJ5k//UV7w/Ukjms65c+b3
QxwZk7MTsUyh66EAWUDg8lJUnLeYtEDQGKrohOp3X/l5vFVF09pGMXi1ZC9Qnf6VkpIJu46LnYyT
892B61yegenavan3v3MCEYNoqC8u/FlhrOwZLaKiZbTBmZQvuBPaiZSFvQ9jU0jUnni9nJy+wCX5
/wW/mSvvms/gcpakV3k/zQQF381Z7cqvdR6kpDvEgx2ekYjzRedxeQS5LFgHfjxuFF6tSezP9/qu
OI0FaW62oevoGU5dTcvD2hntZsj482Je2AZJKzAeYDo4gbnFTkV0I3989rE4uYLh2kKAkQrMoZ6P
mqxrrKzPTjaTxLueCvKLMT1e2Fa4wvVldPuDhJxz+GvZlUTc7F/j4nWkzQCGLxL1B/WxuHUl3RnQ
khFs16fqtTC2lkNqGcSekG/HKOO++7e/g4Y2Yr/VYHItXlsWkh8ntC4zNAZo/7wtyFLgnjXBZHq7
rIS9Sy0P9Z4yc3SrNBg835zlGjJn7GD/4BnXZrTZ8/4KnNa7ahrIidwf4+yolDhuxFO7Yt9JEINI
+fQW23PG54xBwI83IjOBdOL6wvVecjxV7nE7OJadOZ729Y/LS444kHI1Vtw7WZmIYkfwUfzLWCzV
GGx9fre3z1sDepJeOaEUHnHvdPteN0HF1UObflndy5cwQJutARB8g3n8E3ysmt81iQ1kP99wWsRL
eT+zHFW6KJtkA9QcjxSy4grRPeJeiKKePsh/CwJ1lS4Q+bJdIb+XFV8FULtUQUlwIBrn+Xvgr2tc
sQB90b9huN/yw/lPmvPGeFEfsn8yELJ50X4SDqQ+70mcbKlwvJAhDFAUJ0fHYejqQI4FBdQOqsyd
Rn08qSDVL/OmurvHCatbN6pyvD49bnQIKYe9Ue0h7p3u9ScOjMKAg4ZLiNvcC2KoZPgPojTQzV3O
Js8401dvp/MqtqasfsmfvmfECxIhS+p380CLvLCl2oSN58bK1GLk797opXL3k+5anRKubz4CS8D/
oDAPIWXeo1Jrzhs/UuqIjAjgIdC2nDdRm7IxVrdtNO6ztEjpgwMPUnKqZ4kIRgL4Vcr6IcGywErK
Hi/K+g1eaEZFIluC65ojd0ZGiTdml6G/1Z0O0mNWEaMHgq/Bhwg7nrtVlCucMRnqTZm/N7rjX1gJ
ayx5WxRah8vKZbXmcNYkrhmT+30KngWolkO+gQIqbZlYPtsM/8BfgUVL9h3cWaDPd1bSkg3JlRqs
O7NRCfUDKrGFtk4XY8fzV6Oz9FM64iD8N+wIPs42mDP1PF3UmQPbJESPb33qxnv9ApcHIpAeYV3C
8GWGiLiWvjaWs0clyvIt8gM/jP+kL7saDwx2xsPlRUUir4kadYrRoLBRryi8Hncus+xPbtsVJteL
IdXtgb93RHIQXKvKqNgDIJRpg64p9In/hOPg38A/Afe3PS8Kl/DcF8Z76/EtLvsxJx+lWlqsmdu6
xLbaeLPFTLDjsmjoSXUK10SmP8GDdD/BDV0DhPo/EFniAGS3H4h1S8a49gbY1zO32dFEZmua4Krx
nyMumcer40py/19pyV4z6bO9Sajt8vKvcUN6Hg+EVEwY0es8X2m5s9OLARCPpecnmj3D8vrUYPeE
iM5xDUnPMkBZm7f2tJLJL8Emv2Gh3fcc7gawvJSkXro1ajI0WPNuc4fc5Wjwc+qM24AI3DvHFIJy
Kvyo0rQ+pyy8/e6PnC9YRpz9odsFGo7Ds/myQgAx39smbOynLmDtCoHwVjVzeREsaLqwcc4LRfGC
40c/fUK7tMvfsOCkcqk3bMu8KlLMH1/BjXoISZQ3X3A0zrm8aL2dSzYJ+xmuWBAnBfOD9kGFM/7x
Jxj9bHS98sK/VvlquGticIvn7dPgTgrAngaUn5LzD/7leDIKhjUz4YIFaZ52HKnOoIujwjqtACpb
5x3OxA0KBeZ+kxia/T9scfZC3i5CtT/dnxdeiSXPXelmoWpA1LMuaProEoCFzkS3G/Cmnzf02L4J
cQRHwRE0/LiYs8sjt7yF30E3pDTPA2H797DM6ajgcl1w4b4xA9KNkvbd8ayEz5V7r7V8jXQx7vwa
7fd4SYBy5XOZZsKmbN4hm2mqmWDZvNOUPQlWD8RBp4VkXJkfVnUaYMnJtXrYWR3ZZiooNxebWPS7
ysUOiR/t5uwrFDLXDWl6hXxLL6jD01z7J5Ab7aVK69HPhSq5xe1eWBJZ6eQbqukHngNawbHyxnBJ
bW3hB9h80RUAAwg5WQZY0AaYDmAizginN/zzHy7Qkun6Q6847x5Gz1uU+uuo7Qquy5ZU7awLvc4Z
XbwCL7IjxIrQTWVzYIrYCUMd3fGrihE0VosQBuLVxHyt9slZZtlW9QoxF85kSrZJeHPVHTDr+/xJ
3CdBIzV5iEhUDqmJfMCxrTknxaeugi0AeCPwGdDp6WSOAObVq1tEVtnwOwReKJgWoMa2IXbXW4gT
KC/plpOLHv6kKnvivHFBD0Dfbd0gCx2yBeOcPvBvf4vZwyVsSvUe9KTJ6eeyYoK6MDj/kF8lgH5G
TYDKFLuJhHbKVGRxh0Zchllrtuec26+TiqVClNfec4SmJrTdR43g+RPOc8AaaugM+ssud9vko3ko
4T4WLt9SZibN2yhIrFZ3+adQio17/Fw9phn0AhK+ULI0iOsNSPnF+F+111vtRjTctsuugoLtBS4n
khCLZ1VfbCbgeTQLwldS31xHI5auqb04e1Yc28HpO/T4ncSXzFKSD9RMKjNkigWEY4NiDFVgllwu
D61MKD9HiMLKIjtBX9dgVLhsJHY6YJ+l/B9EJUYFNPqsUHoHsPldy5U0Fl5b7Hl8eueZvC5VKa8d
J3MOwDwqy1F3DqTI4L3nQN6diScnYj/9bUnNQ2/HFYy41Q8pyVFD6b9Mcu+V59Od4H0B+p4ve3rE
IG72r6H2U8RYwXgnqqdkjrpNZgkDbl2mR2TfRjTcNK0qjMM6B7tiAd5CLdpR4OEfmRpGFX/Neygt
3ymZD/o1g58j8bhHKulKb2+IdbmQ933tQppgbqFD54f40ebNE2nVdwTUUyCI48DE2Xd4F4Gd6o0j
Rvdn6e5uLOywZBmp4L9Yx4Kf2kXXrZPg5gB2LGq5RPckDrE+6Jo1YwTozMpymGp0SRlKDe09ulZV
TmRI+3U4or9d470AV6//RhKn1bRqZawAIFM6Wn0tEfDK81ludq4OFbP7uVQF0BUpaigeqEsVA1Dh
Qt84ieDZVcNNP+7Fa3IFtz9ZKB7N0AGQqlyayBpP7bZfe7VyAo4awDCdhIv4ciDOObUpBxSIZUl+
MDCA9BbRdgqzHz4u6uoaDWOmN2LGyKyMLi3PMDLOsNc8DTJZ5wT9LAATWGmb+2U6b4F2vjUk3txk
Uz+v/QZrd+iW0S0tS+dko22f0K5TC4JRU2TkEoBdjkxoztACb70Di6jzDQsWFWrhkvVGuK898vdD
/47rGwHw9gTe8aKLlM0cfIOXgRBIRJsTAKnz9qK2GWJ1DwTqWAqUHDmPlig9wcDHe5ZIVeaf6i0Z
lCKyDiX/zcDKaq3jXg4fWz51CPMJUuIMP5de2f9pV3IsEtbbKmwMKkdZ1yX49C8p0cYlQf1sISC2
q5xlNgVHA/MydOdXSxAHml42RrLi9Sv1wgY2r4EGfgdoF7KiGulPLqpz79Xnwl9VC9+iDuxkxbj4
7OywNEacGD7NbhO7nQa34/j0k8qVIUsIlV5JSZkXF+mm+DccOYEvAoJVU0z3NicDYvFPLJ4gaAlx
uOyWwKT1HXvOExOqAa+c3bc3bPXPotgIKYdhSCITBxWqVS0UgxrpcYe9Kh6YikF++jPnho3+NfTT
eAWwqjjOvd0KJb9jFpdq3UnYblpKCU7jewuOQeaPi9UvDPs6yjJiYI5E+wnhrO3Ie4ty81MQRFY6
sM3IX9XtlXp0gl71MbWQQKUlEPEQiFCI6qHTYXvwhrhTQgPXADnVi/TlzPOzfn2xiJIJc1wCSilo
neUwd8bat/qdLL1XrBaDOIWIWSt2UquynkSYxnEwVRh4mWMd3gHm4dtLMgxWwBh+r+mTpI8HjG0R
A/EhGBkDlDv/MlFOK9IKuEcDR6JBSLJkeekJrlslt/x7aqYV6UhB9npvN2Msm6XjfipDEtzi1YfH
7/CA5Kx4LYlisgObher8G37YtEQJ4Nt1KULesJcwsnn5hC4Y9LhYftItksmvvq5XWd0qs9G3GH+9
vCxEhfqrSwrmcIdVBqckgtBs7ziSLQe/YC4lmAXkIgQDnv0xb5ru15gE5NNj6HJQ+kdXZlYWGhpJ
abfiD9KjMNKnySVuVuz9oawAfqQ0RoVzhBijG3AZ5EcQDXwYkGSCTWCOE3zhhzwDK9jUSEimWXIM
BYOU2Rw2aVz75mCWrw5DKBRHURANb9PkZuDzyIroFkXdRB1hP+xsxunDg/oiuAQW+SaN8c7dzZ9n
DLkFA381ZDu94re5k2oJ2SfA00oibvcSkYSTjUcnWXnuVctr/YHvHY92nJVMSFsI4yVPFmXCKoxu
AYQBvUAL2hjfdLgyL/Ys6aVIvxq4yhNa2yzmlY1C7I3dr/gJEwR+oG6Rntqzsob8dOuANeHuDv2+
UzLcx3HsFW8knyb7Pw/WBs5V6bNsrMvLZIIQ00sNBUdEdgaipedmFZUmbZaSoWallV1Cs7X0037T
0I9uPfm9d29Wj1HoEO/xDJdZpXKzsghjZVXlSUxPUvL8RuRDO/9BsAHwutfBEeynfK3gFQoYLx7s
HC9hFqmOqy/9shgjboKgF2/zdVyBIH3RMSBW1LOSd51wzzldCUpeH1163Z21e01aSuNfcvPYcm3c
9D4hgHy/ZPqs7jgZavWUNIlltyFEl+aUxZevYgvRcmRH815sZM2VW+dJdd47mwBkRXgwAUGp1hCH
ORBLPT0xaJ59JZk3DrtNB4ySGZrpwiwr8ndK+UBR1sBxX9asXOF+7bWRN6+wj1GvwoYQMPBN+jmI
otXK6Gv9tiUd8cIqs+pT1hbI8RaBtRegnWEuN4dAuLslTy1AvxkhWBE/VGLqYaTm5iASqliQ0VpL
C4k8qPTOpWFtPC6j7bbVnElEJPVgxrgtcjck84eMlDNQN8L7bH3kWojdPK7tt5ut5ztX1CVeDbVY
uTU1nSOlEb6f9eqoWAtE15YUwmYNdJqzohadGw7vw0AOpC9+rR85t8YLMG5sZQsZP6l11ZcXjrSA
LlU4C9VL5KotwN7VfYE2xUTDzjo9fftwqZF1RelRpdvaq+CIcSExdoUuL1UZSRJxIbqoGvg9rm1o
z8FbKR1b4r4nYmkqIBlaOpDwp6W3r8r/vJvHOXmOKmrinXUIwKzP2qeKwmv3VlFVs8zEaOHp1TRY
ZOOoBih1bKrUh2M3TGDxrhSPjIQ55kzxnluWy5sXPIzcLap/duIShrz4LrIbqtG74bExba9bi9LV
LUyRmwvZE3SykfSDbaTiw6bEmQCTLHZhwa+0CgH+H5u4rs9hK0uqayEN9gCNxnaqtR8SC9hnyUTM
AEmrNy+vFi/M1q3H+ocxyzkkVt0whjoQyqRNqTdHhZYsD3/jSza8AlMKB3g7hPGytQT4fb2dWDr1
JBpZudXSwMiog7Mj4kezyK5q4HO6U0DrWPjBqy+5luvHbQoO2Rw4gqIBhUhpkodKGZIb6Dl1F2uA
Hkh94TW94G5LhU9WWwROkDNLlmOcxfvnGE3lHFebU97uIQTSti7t49XZbC4tpVgQIR9Cn5WdOT/h
mX51KK1olUd3QoUAamEk8BEO2J5EVS3CT2KNKD3XtFdxaqsqctno62I4tNH+MFN/VSGUrjWiHzzB
dgEYn5aq6lec3c1S0kwUoAdZ1OR6V2AtDS4jqkOIltkFLgPLLtH25GqjJULHIBVCnjbqx48cCeBf
8o29Ca7xRP5u/b0vEqy7GkEULTPRftf1N+qrGf1AOSB4XtCvAKC9/NBsaTGCkaK5l+vb/nqli7+Y
4hq3wwtLePRjNXTgFV3fYmr0x8R48LWnP1xhRyPbNsKSTyemUb6QH2B6PuZ6/FxOu4P2SFUXAU7J
WEPB4ojx8lPNn/YjJEQ8a4kwr8kX6h7WXDkIZiCvC/Hu2kPYa1RFj5eUF6Pzsj6dhhEjgY1JwACR
XqoOjTRxfV75iMyclx857wOHkEh3lOng58rRuOGLrp44Ty7LZFBA85C4qQWrIZsw5GVaufRu4tDJ
ZYKblzhUTH2INsaKgUKErd6eNq4Nnze7hHDjf3Wj9r01wQ6WpLO859+I+a3WSGUzIawSismCvMfh
ZiY7ngpaxsNza0gHUTK2/CaOlYBUNL6H0xLrdSLURrdCkWln4ZkJ7rLo7SHp46Y7TRNgoKY1Z7z9
UL0WklBaYkhpxa78Gg80ZR0JpXerUjQJhY7K6aTV4st0CpA5Gn0gKlMaZsktrPKFMqcFMOPWxrws
krNp4mkVdjFERoRSJ2XqN8PiHr1bGpjlBaNA/99Tqr4vIpkTPOjUOesPwAqo6hQ9GRl7ARXC09QO
OkokoT4Gd9/qPQWfJgQsfkScN7UanJ/N6FN8YwlOT/ymbabLn4/o5wowc5l5vkNTmBAFi9qCa4Pr
n4i0Ddzg3Wepe/USIlfx4Tt0DTmO1FekhDwpEF1EsL19iCz96YYeueuj+9Mb3MZYf9mHwn289ehX
0eNKnkVtdFU1ajnwX1K2uON05Xx/P4UY3IMoQcZANOnYqQUeASuvKldyLHh8mnU291BWAVI+Pm5x
3eSVokvzC0YVTDm7NFgSO+Ih7+SIp4c/8WNBqZWRQ4pXWj8qJ7vOg6Cfkh8Y9/GKFLtt1rlw55/B
q0Gsa+h04UvzNxODfcjbA6akgo/9E80ulDnGdigT6+7iX9LkW7eA5uYG8b0zjUcts+r1SXTGEs1/
Af3T7iJAENHExzQEgFHVo01rHtyu87ebmyjFCzt2SWHwkoQEdiOS59YsKYy70ag6WgfDLV//R3Ii
6ly1hP306TG6ws2TSBpzHx1ahzRHUr7ruUYSJvf3yVCkWVvqIBchO15d0WROGrglh2eAGP52oZr/
MRMQeO4MwQ7RPLWoZYCshHaylduhnImxlFAc8SlowwcjASWerSy9+yLZxuo89UilNO/haGfffzvj
VJbYPE6f+BvyUanA6lIektomyDB7+8iXNImxADS72TxnMTjHJSju1saeWCSq8T83Se2XZMrIEg06
CS9abTO+LZwkxWwlvFqEumDNxVp/Y7+eDyV9UwzdBrGnsqkLRKdABich1pXcXr7MzvxsNnVkFN1z
76DPzsquPJJ5EVlihx1wP7ah/Q0WSA/5xyFTimCUDBtOHJLjAHAf2Eiulgga+0xKwSdNJukjpNX1
/c+HnPupYSPlWz/3kpo85d5HhmJKVIaP8zYlTbS7uRiVNemFyXQwyw5l6OpWCfOK068zcKP2pPtT
SUThAyed+kC2lWzFziz/u42dG3lkzKzqhGeSSZdcVTcD6jM9PYFlNe0MC0eV+IH6Dokf1k7qliFg
11sxJgaz1Ua16A3BQoscW/RIO6kCAXCkWMF38pxfPWwmpi+8b6K4eYYe+TgObYNh0ldXiBJmQAfi
o+9/Q+84Xg674yzHcXEnk4G7dPyxeD26vspou9XNIFl04QTjD5IxV6/Fr6bIvxcHhmbT6t7K14+9
bidM89TOEAVKHgnk8pGa4qV6WL7U6f9k/DMWXYWPDx2bQ1iuldltfhYpZLlvf5eG6xibBy0q6/jD
uOCrqbNMquskRZY/7HtBdZdYd7+mFMpxddDIx4QOSxJbZcr7b/SNr5gJRCr6/pr0NIw9uKb04avw
orESkeDNsiUB7r/kUjX5ZmOuoWqf+7fr8drlBirIiXzMC/l1V3eahw9/ez/xVm108FtGgtfIXEUJ
z6nEpeTw1wqQPgh6lfKLBYx6Kv8ic5IXKyuNjdpyePdCJo3feMBZJX4wuAQYcoqJLzLAQBaOn5qV
yGo+P4gcrl1rlURRRAOsbn9VWYF0grv/BA21KL7L8NFenQLc2SO2mW9L6mjzK7DL46SNa67raeJx
lCNfuT9BL2fLLEO0N8An/3EOXDEjPLfuMbcFGO+N4NKhxrZVzEJsTWBdxZd223olIwpAj0p1M0X2
L9gUhjyoV+03NlB4CNWLWoJGlAis/M5d3G2HT7qYM97+a/2rKjjvf7Cm7eIaYO+jLWngdW0lggLA
aM4TU3E3g9pqln0p5Mzvop2Bq+r4Aco+ygmHC+v/g2Ok8LivjfFXu0ZWCc2wsOQFCmcb43FjTvCb
KZ6yPPPdtKGDPYT+RZvZcFRfG4PN9Nf96KtV2TqKSy3w2g18edMOjCH1qhfocLBA9o2uNPCs/g02
uRyksp4jbzCnE00OoD4MQ4kx6lNAmmka/jFxWcLw2xmXhVCrWEl/gbyTDc+XdtjirUa/d6aNZ3o7
7Tl/dOHc2qhIy93Q4S8mauJ2o8EvXbd3GlCRAStL1kP39Go2BDbfOLljsiOFmegzXMhW8ft1i/T5
52Hgimbq0p+PAjU5BbHW+bo4CYITfwQHCq3dchUxlMxDCWBsR73HNb1YHdhxhjNuefoO9vQ9duDP
5x7vuSJMxxTF82OhefpB4cl/s9peHEgWgSwgioD5NipH6Q1B7LhY0toou6vvBnnapCLTm7C8FmLK
WuCkoTILyPWELcrAAFzfKykmfl+8u3o5uEtn8Z5TrrcFZ/kXHrWHzBFsBM3ZsZCPT/Cn67fuqa1j
EcTyNyv/eLyzAA607N1V+W8bVpsZe2NrrlP7gYQG6AynxtvzMrVMrGvtvrh+ZFiT2waG0HMlcH8h
aR7JY+L+eP601sgzjeUzv1cW8KlyeoqYXpRuueY7SV2EEFPJsK3ITQ27PB9lA0vo/tbIl16pgKD5
dszz0gty2rwVxMLfDcEZUYp7i3hcr+qDSCFk1m7+wDvC/1QDk5nxcKjtKYMRc8aEmutuv1/iQ23t
hDLFBqKuMLRRiS9FzKffAoZayAtBC2biaYeK5ccqUnBICIYN62byf1dDpWX1C8zPDnFPYJD7S9NW
BExzI33ZHCwM6ofLpJOFM2B0gnQ2xK8bbvdOzpZsxlpQAKUXIoMhSz0N5sOqjMSbFt7UYWjk8dHY
lW4gh9hqGbFlRIZjEU/WYei9/IENKojx7atKhp2OmrFmBLbRCH6efQv4y+tEYd7wP1PRXEHKHdRm
II/B0oNqmx5p7/5cYJn2u24wNQ9uV9gsdJwnxTTcE69WaZBdlRk6JM8Xn6nKMZ5ipQNytCxgSi6P
7LQen6bl4nzLIPK6iYB5wTrhBmt3b8FMzKnxf2LFDKpSuXkJ7Va2hU4HHy4fzRWJ7HLqswacD1Zq
UROazElUBbizjvLvlvIa921xDKtDc5E/OIJDa1w8yTIr/SbB0wP6Hx+y0Nako260KpmihVyeAiYd
nQqiEgVftE6nSO5iycZ9yHPs5nTkUgfDq0oG/Poq6/Q2aZzotWlyAVNLnBtK8W0CjqQnX1LQX6xf
NMGep9O4vlTrth6ohJUmPssHASoqpiNHYgbAG4NDgyqk8XkcFRgn/kcM8SIMwfpSefqTUXPq9l37
nRIdu3laJKbi5jYcyvgXeLuFiVkK+KW2UFQLXzYI9Cdh0FmGDLr6HmdMTnvw4v30xKqfrHRWPtNm
5oTLfGYjz1bHjx5IoXttG1SLjsQ2j550WSCLCagPjyj5gDI5CbOJq7Yb2+8SphhX5GsfhlOtR5NF
//65EznMuPeX2yWAkmQE6LNyg6XRQUM7NX7HMopJ9Jx2ep38HsCbtdQdNSUFzWXa/ZBv9ByDAmst
VQqjqypOmF/AqJfKqqQ/Lo3OppiOLPkKE0xxDsPPoreDmHNumnOr5US1h67Ce9Xh1auymiC+T4TQ
9eqW/v5h8s7RdY2VniAoAycbE2LDzhSfz42bgMyIbIWg0H9rdN7Ylf8sMK24x6jEF/uMOwpxg3f1
HTgWnya8AHaWjBjbqOcBkvLodcV3IGgMsiKcbKXa1Czo2osk5rj4rLIaoQ57dRvMlli3mfjCZHrv
yrRQihinugAPXFysUxeRVOW4+K706+dhr6/06UrUvTsyz6rOZ0F1riP7UxJzO4n0c39hFCEdiKu5
OVOFKxBnw2M76b5YaW/SR72bVyKp6KLTit/f0RsytNweT2+6d1PJcRjfLZDYcj8AiKxE+cOujqtI
gJzGJJo/3Kln6aQyAwSdTHLkmZ8RoAl20BNx4mqOk7fQTZ4kufUFq+Firu5S5r2vPypKiWTBVZOy
+6sCWV/7l34oaPzuSKteXoh7HtDl953XL92Y3NZY7/zNS789/PgiXMto9aEIQtrPnwOW0rT5D/WJ
bnhHKA75jXsMoaJVyZBgKY1pbH6z0NuNk7zQA3jFcI2IEydIeNCBDqEpYQ1ecsxmuOI9kDz9QP6l
SvY/Ei/iOucCHkgI3OHwbRN0JgI398f146pQm8sfsAxa28lBZVB96GSASigWtpri7HwyokHqnUPI
OnYSTbyDskp4E53RD2IE4kpBIeX962WzgtL41WUQxubZvC5/OPEHP6lyML2OhQVVVHCXLa8HUp0z
gjmwpAiyq6ci/hblvQ2gwDTdju3lgir2dnARn7XmOlNCkuV5Zn57rvuXZ0HfGAaSjTyEFH9+gqu6
opTK2hIEhsznc23Q94WsmeG03iSYsNjeqAgU0rEYUpMhyHWOUzKmtJhk7FAfsrMkTihiTdH0yDEm
qEVmvWihCTUTdEQW6EALNtjMtuJlOy8LK408i0ov3cedkcHGCF6MQokLWX9cHG7nB/4UzHlScENt
F9oPlqrgc231MUDuG8p/R8bhDe5Zv2NjNDZ9mqG9WJQUnWpH15AbvLxtlWwHwbFg/LIObVMKoJ6N
k3f3VCuW3jXdQ9dxvbkx3zZXHJXqsoLXXAV82d4ocw4T3uQ1RIe6czA7mY9PyV8s1YxvcaoBJTS2
MkMUKcqAC4tXBk3nbGiyoryX0fUzFkQi7d5U/Lsj9FcamHNgb2MgdrVRK0qmtftyaOgYDm5tKMtX
U9PO4P+ODULmfoCrBLC9crX9DIQ0WIn3jtWpe4TTCXWDK0RLSSiHH2Tt3Pn691Hb6/KTOwSW8sCp
IK5PxKyL0cVOa0611yb9RV5BGoKcPE+YiFBVJBoVJ9oLJe4ZlSQroNVh7hYHbBAkXzJ2R/p33Zij
thkdv6zzQOcZzTkbs7leV/l/WNjVsB4uq6MdiFDFgZkthK1uzdWjbhB17qRMwbTOKs3+JseCPh2/
R3zKxTNLg4yMt4tK6ClDzAoIO2774w2WCo+5eANZWn5Fcm952vdVKv78x6B7cne2nUPPD6aiFGk8
ePJdCYWXpNZRpbILYrsr2Wjvsc82aunTyB6TfQTWBIF9826LzUGitLdnIVtoC4BhW0eskisy3WDq
p4d+l3qyW0oK8lIZJp1p/zWjLC1K5CsxmL8tXmL8wFpg5swFb85s4u+8402ZUzyANW1JLkJSluKZ
OvkckE25sqrSsLwytfS15MaM+9hQqWXNopUnmj5tgSb5OrYxggcmJ55PJtHliTFleK0puxP9ybBt
zltKzh1R/B/PAkBncX+hp+CzbbddpSTNiykZlYpie9UszM0nH0tXKQisaoaYUQzpCFDHhnJx8QtE
yAXt+MDrhrR11XWmXmDJrYhJi1S5vh0wvV+9bqWJBjFRMko1BTlo7z8RzM4JylKP8QwmiiByZ7QX
Cpeeqj1YBdpfQ+N9IjD4jQKPkHVeo8ZihN3jEeMsv2AC5Tfz7nbt2vxdQyM5W+kkWqzivmuycCnF
i/D+Z+Ncalb//h46pk6OpropUM1lLiQFXyHae2CYbhdD1nJdWf86RVJzbgKy8QJtT3jQk1qiwTMG
MB8a9YFBvSKWBMaXXnsxyj5UF14wX9yjnKnfqVkkKzxfKuSsSSRoOROymTdSe/AptmCy/7RT1f9B
zKuH4flcHZGUeqHoUJnVRIFXGhiB3uJsEaobswbY43AjGoD7m8G+qcFBW3qGbc+8Z0X4GogZsaAZ
4rucDuE5j+bMWoIkiaUDiN20aMtB6ZXd+fu5nHEFXSqRXJHiSZsFowez+KNUI89ydo0z89Ja26hT
aS4RlGeu9ATV6yKuSRJXFGgwSCBDfBhOs057wtjKfOWTNnjFmBRoWi6AJd4Fcg+rWxCqXZ5s7dx4
A2OZpaQLIolLu53RETxifWZ1YxNtlDX3/ojUSwXglDMFeYQFLj27ox5PeqKvR6HU+ZKIwn55zw7u
RoeFK31wW183x9qyA8MBWfzCY6rBfiVhaNNFbvIn52eV5AZrVk5Rw8xXTKFv8f1dmGFU9cIJJisu
Yr44cHAa7zfm6hwUdSaOqQ2wWfKPMJJZnwwAVEzlXTA127JbJEZNJO/Il7ZAH0i4m6rQ87qehSe/
D6rChojHeEnXqPQJA7onM4YEMY7N+7d/qs7WEwpxs9VOYhYMyMGtUEMxDBy9vn1/x9DvhVt1ZNVi
v5MEnbZswXvDMl57p02yyBEzbthO06tA6nAAjm889atjWoRyQ3ZAbakaXgT6NxjVoq0CRL72YOFi
KXKDfx8QNqu5CZyGepMp6AcA1DRzdk2xzMuKsVJlbHQv1KPXCccqj26mghwFOmUcZl7W5twM1A1D
JNd789tfkIgW00bT3M5XrQYe+DD1bH6VOkJdm/yF/55MEwepAOu7WkrRUVP3I5uuunhkjikRiFNl
l7bwtxO+pm1Qb3F9VLL019nFo1c5MsNXPAgvqB5BV4vO7wFvrgpastGW09DBvRV6ruDMjtdx1axD
6hhmCUpf8Sa3tmVcGCjS2p2rVxVs7+iDIJHUo/SuSft2jeBYsyopxgu5jajMonLfCEu4jZvA0ahL
GmfezTEMeqYZuAG/Y4N+mGKEisqwOK0kCBvlt+/qeLxRzD6OqUFDvEl9BkapM1BS6xzBh3SS7A+6
9RxlK0Xsext/xllJEdS1g+tkXU5R8JvdW7VkdGApb+6N9H/n5Y3JCwbFA5yS//kntbjl0sjU5TmM
i3KkHabM6X6eftWqJbvcqx93YIp9UnO9kJvivDS1fmOXaZmBB+O38B8Cvw/e9j4aV2etFFO+WvKZ
rhboEP/CgAsXvKjv6BsiaD7Wqhh0v1ZVaR2AuptowasmybOo8QYRYsnHrXci/Fw10Ycczi8wxgVS
yabo79+J4EADH6THp9fPHkF+EFwPxJTojLdqYYa0rqptqbJxbgPSFYEV7m4LnCZ5C/u86l59fKGb
co9FZGDVA3dFUx4loLENYkImC+Xq2+5MiDwHE7b0w6IJ0EtxdVd+aizZ27dzLv+qqE+OZmOoYxd5
iaXWn3Up+uJ7OYuc0vXq/l/HpW5KbKmBjT/RtIC7yThVURGUXfpOWeholIxRR+otPkBT/EhGrwHM
XmFC1m9zq9WEZlJWZTLlYFxmClaD+eDIWVc2kuG9BuvYAUDreNVDUahBZVuILJloSHEiBLThqqr8
PSePPWKdDs8DYKqlFmfCb3qbkN26hMnhHcmaZNJjssIxvFPl7rNK34Sbj81L/qyPDXHWUHRTP4AY
KVcIdeQ+TAr6UeHogicI+ca2neluQVfq9MDA03emuKVSABre4ABxRUkAzF3Fb4CuegAgRvmRgm9p
+iZKamjgwW+lX0sAHG2jw79ksQkTyM4+hcoAZuM7CWhHpoIkADWmZcQAzKx+PF8y7Lm43wlXIyn1
knUX/B0sg9quJDEexwit5tvbwBdZIJRwaoKRjiOzxEmTxM+Q76JBvaMXi/kbLEg6LJwE3/vE5gNG
dhC1YHdarnpFs77aDcsnkiFTUJNnEfITlTWBlNPpyWbVwDZpJJplLmYC8DFOD362XxSqKq7dhN7t
UoyMnbqVFchdiWUTiChWgkxl3UfmYq3TU56e8Og/1ye+Ab+5HcFEGi7NUihyQgVmYtGLk2sbSGOW
p2x6fcacJ6K3+gQYr3pbvik+rgTxv1LbCRBo9cJv/w7Jdq2rvsqfpwHbMKg++J5si/vLxEDzBBFe
sjtQfPRdc7xaSGiCo6P3HXBeIXS2H64/nsXEUB6OHjULero+4HWrNdiXZPIp6JZ7oAfHZT9gT2n4
y9nn/dQuVIWTWT5UFAKg6Lvck3L2uwHY/vls1+Zeaol3qQIoCZL2nNZG6QjBJlZ/EKoObBCsuawr
/o5w3vPPPKV18Y7WA67YJnBZGhdajOTIDUu/CCOjkVvSBHcWmUGTjT7FAuLfb718N8iM7o4RmjvL
iH33n760SBUJniXjQie/wmMwCbpUuJxnJgI7lGVG54d2DpbIOOmLqqAp0c6A43RZxZZ/BZ/TetC+
0rMrkVfjHu58dUWd4FDRcr6CEPic7kQfCJzDB9eq55XzP9wLFXMV3qqBuGNdrvLPJEok6IytoJZ0
C2zqcJouNtMLKPi9UG2PxOg6u+MAzYHz6Dmy5isD/DSQi3BlffdHB1wJ/A6ncZJsRMjkdmmK8XMh
HFk44CWEIECWygJb8e0nZrfyMzc23yk5zZEjydqAHHGdsaQKeKTZLci1wbMjYQxM+ifXexlKuzLZ
KoIVSbEzTXWIZuQPlSax1au18h7wvMtq/qXJ3VI01RTGSJzalUXhzSOOMf54s2lQU2DLtJnmexld
0Q5tvOGuzcRj9bLZj2QCzPK9pXA4/+b50oF6Ig9S4hDjOua4JKuwwx2pq5QaRZkNEXEo6jWB8nV8
oGHBgytndXgE5Qaw37EZxAClGC+95w3ljlIPxnTVMZi9IsrIxl+4IVhRgsv9eXI74nzeHrOZei2V
aCn8m/1g7xcgLUmqgHFpZPRUkyuwbcUxTqsjHJbSPLmEFcSlxsijlvpj3GXH2nmHOGKm3W+nVj1L
VIHDK6bNns4IVyfAbi+2OgNXV/6hzvUkgPdUlfNQMFAnJ0AxUTTxxi26+VPCGTFOkNTfB7N8rT0b
mK9a3R/yAd1NjbnwO4KIIKSsKACEZ/PDbTV+5vjByJgZJOXPwji+A3zqU7ybmGz2i9oQimkWmLe1
A2Z2ZFXZu4EHu70WP6lE5GOvIlzZYCrgIuucL+LzpCSJKr89e3dgNm60smvULNTMgjuF80Z3sk0E
Papntm2rzBXu9AMyMPESJbSJd54jjxpsmgNlCF/T6h4CR0mjVfrx5xDRg2VKh+5FpE1C48uoGQWB
1sA51oFnTuBmMtJHdor+OVmW5IRSy5C0FICflWNUnyLAmoSKXJ8RONn1CIS+yTUvkrkCi54lEvkg
weWG6NSyCqiBPclrTJHdVQ4Kjuf5h1ucEOT+7Q/DC/2amDjfDhRb/8s4MUo0hE0RWkBHoCkEYwVl
gtlaaOyr1KVfjM9l69MCkDGAxpzztRWhuWo+d9HMiE5GfrGPZKFAs7/+xbks5jPnKkrpUAts2vIZ
4c5w0wWgXuy+F+50ovSIxPuFtpG97hzoaF3Bj8AqDzJKgaeDUEY8x5QhlQHLv+X3ZSHRZEnfbjM7
EW5YohkCF3X0C1Dt/rTBBy6hhCV26u2De+Wzyl9aC0pfwvNZEyrXtkMHW5qS+GjK1ph6e0I7EQ7v
nmGw7h8MfHR8SrbhACO/mb3I4sddeBoTK0wlRVng244ks4k4KgrwIykhytcIB5v0VuDZrl4RLn9j
7p6rmx5DLNWKjeXDbN+pDTVUScuKbXGjLEkHbcWnuNUS4jCG8grGnQur/qT7kdol/3E41jvGceKp
h4hQXZE5Wvx4uL27J9Va4Aw6d8nxlLVwYW7MVyR6bY5zFa+/b4Tjp/spQIKutd3ERVMZqrJh/iBh
ECof2psi9qiik2ZBtmKYF0ZcTHgA0PlWi/8ejrOF1PW5xIwSHWfG02XIcwi3ju+JJgtWm/e7vdqJ
E8yl+VhULCyiUgWdAEXFSBaGN6kigKynTvQXBiAscVk4zFpV2LrcksiZV1FqMZrZZ3Ohk4qg8n3z
T7sGkVBAgPNuRjAKNoGw2qiA6KOE5OyFDQ++sPNY2uYUPrX4CGubzqrzglduUx7gu0FB11F3vg7b
UjY7m8u+KyCZr+rwTdY27IeUuWCB+K6QHfvDYMos47769IUN9exIkQ2wS2x0LGtyEneBr4BAW4BK
qfAA+1vFB49QNUw6zWOj4ByecwKVdNIALLrMq/0Z+EWqfoTzO3HfutqFB8DBrPCLJoIznOXSx0tG
dQm3NWYjvSIsaxC67cil5JUXvaFageL2LR45HOqqf10bzevXNgYBB/H86LQeZdLmHPm9B2QUN1wP
NBZgTOzHfWqZpue8pZv2LkWAQF5ihsEtZ644NOaqmt9KiF5XPmNJKAexwkRfV6ddU6BgZlID5OIw
ZF7YtaEcOIzFj7D2J/7xHsGkXzGtfqNwurs18vFCueTPFlYfmkdn1wHLJgwqw8M6fLrASjHfR4wx
XPAS8yjWlxOfdY+a7sPtpZCtrSQylVYanrVVA1evYN+Om0ICixOv0rQznMJFczMFya4GwAW9bYgG
OMVUAHQ9UKT9QTkwop8SpvO+9cuAIIDntI+o6TzXoyelShxPgJFDA2MqYoShhSFdQWPL0sLSGGxi
yUw1aQAPHQCqktWGSrjw8vrNBuxgMkxKNDTPFQNjwY2z9yf0w6o03YO325aCpJqBDX8QtW5JJKqM
xZJEsHrVVj0Yt0/RT4vf7tDGQgjPggrKLRFGQ5OeqhuqzeZXEwOZ2BTxqoAumV4N+onih4PyGCpZ
G14T75SybbiUWLx4YLnJsvFOGLGlrnHkNzjIuDU0RUyvnK0QpvyMo3G2UpX48T6+5LVz2PhwNhXv
R0UxoahG1H7wr1StPOAoS8c/GLqp5BdemeCqC8CELZidiguHpPG0Q0xkPml2qbHcwX5ekzia9Sip
vspML5eY8jg68jpJS4+XXvDbz+1fG6QJ59Fb2eNSK4PW1qE8P+2vlIDfiqppHvcpU4BVgetecz6S
3CtyWVWNzWtHsq3eeAFtQNz73lA9soN6JLdRc6v5SymTTBexethZZmIcVFkYHyJcJ5cUDCMhmb6f
NHjNOH1oMTY0iDe9+VtMDqdVcfpLaThc3xSnOvZGjAB4aaTDaOkGtMJkGzyV36TOKD8Wh8jYkdJ8
SWnlbOL41GiLwSZfpwpB7i7Ug5c2PUPdp7cKU5MXKXYrywDD4Z7JDWdW9hW2Zkj7lY2d1Irkz/rp
62jNM1813DeqUOIqrfYDJre9L+9C+yvUh5LXW4eF4aVDXbz2K/XkVFNxcW7zokH2EB4zrkY5GDHl
KsUUhWyU6KB9Jhc+R0MCq5rglDfh/IAXD2ZhOJ2gXZR0hj0bhLQks542HJ9FWPd+5co0lXxi6iRZ
315ufR/MYtQCPC9r/Wd8s5nI7GvglsSBu3oLFc36MElDhwdOt9NpIX6FDkUh6lLxewzfx0cYQgCO
ZMEUnU2HiGAEBpMQb9/fnF+tlsnrAqwXL0J/Q/DcMt/ZF93qcBSmVaTDf52eRySMu+Dkfx1C3GUx
VoG9FZt7tfP7DDBGFotFDHGCp0f8euSnV1RUj3RgvFuptxL8ubRgx3lEyCosAUkl2qAtU74PsRnQ
jqFAaalorpL0u6PtuLhVE2Tzv7n58swCfPhMwuYlDp6b1tBegQedL1zA/ypGZduLxysZb48lPNu6
uw0afN44i/ITySSnHCqDZgQaJVFsqpSfPLUzlMJYAfDSqBlpXIUnZLLapzWoCqnHp1K8RgEYabi/
xKqyqpoqVPUQYmEZXql0myOPcFCqjBRcUT/09XnvGq08i/MEyFFC+HsGX+Imtiy7dIXK1ZpD8g7k
3AM7SnKnCPWYdtpfOds1i/b2e2EmAWKMlyUj4grXTH6Nlk4J1stRJ90nOc623G9qLhy/oX4qosII
OLCNEvNi94zbimUZ059BtTui3HDFRBilEn6L4yFFwZQkB9cTB00CzEpMmw1UUBO5AUqJuX1cwG5M
ELZLh4zLe9RftTm1VpEubF9aVKWk8R/ZJcQHNM7lN/pBz3eScDjM1o21Cj1yrt79ncxzOZRZT+EJ
Kdci8vjmKsIrJm+R3iyNYPAVfLBTU3TmmecEM4Fx6HoaEOIayo6ASUDqafkBRgHRYcIhTvSNNu1d
zNA4U4VEbGaeuXG04ZKledbDN4q22bGJ1usoBv1OMbgqQ9Sfnb3DRkSt6GBROkRQjlAHzCd6eXwf
IFG/YJ+lvbKH1/ikOSNgVbw3uJuGBehqOBjxRZ6Hd0yGXFe1CheC4xIQAyLcGKvDvm0ecxRK60Xo
jICfHOW7S8qD2bnX3Epkub8oYKCORCa/NJhNUpV6J8cF/4dhvFAPAkbSJijVvWCDnsU2z/HJv+ky
43Shj49T5B/zN+KswTPW/tIxLtnyeIrVx+tfxIwYLZyRpE+uzunbhqTcEAHN5mnBDDBiKHwINCAW
m16MtMb7ES2BaGXrYjzI+JieHiAb4u926PczyIfUU3QM2WxeD+XLRdjTrtMhxMljuDxoxP229RwG
3p3JSMdzGpvvcpdAnCKNC5DdZSL6KzOyqRHzQKHu/VBrrY4ieY2aldSWArDHZeu1oNiqS9of704R
TVFjGzSPjXpjj6eRMxCqIgCrUfUucXycO4imWfV8wUsHI63tAKIFIp9KeWHK8ogg9ICsih4cRpVF
WwtHWaqdo+iz56B0fWzSZb4arb9oenlKx662jQWs060S7ahK+nAaACIt9FBS0qJXoSRHNm9ULoki
xcgMblM4eVRzEt8iGelCmZ9SIWoTPvnKZwzNOGj0AokEOvW6cHpcoq8orEoTXTriQXbZjIp47sET
hdsojwZT1QZJxaufP8xVle8zmNn24dZRKE+SU4TXastD1mEYzGU8mcCEjLMSk7NFXOQRTgHQCANW
XOrHTawJ1Qj6DnKsjDLKW2FB6uIhhEYTU/LOHkZMbmjQULVfFkHxGsDY1Dz2Oh/+PJWrTqn3v25P
phVw7VhHruwq0dkYoJQsaYr2Irp0UoJnQrgbGIlD7wmsnsh/dy7zJkVZDU1kMRpFUJTFQGc6YGSZ
CMIU+hD9jG9iVdXvpS1mdNYkxHEGBE2sGadVW9XkppRu/Va/nWOtaMECU4wGTj5MVT+yi0zCWIHX
HHk2Ei2cvaVZWTYUVuOQQZsuTapIqgmY6Fr4J43jpDtLo+2K6XzvqgpUJrrTdW15gZpzFpdWnqok
uJvD/Y0qJjJb4+x2eWPpnyODkdaNLMgclVyjFnrD04hH/HzACg5hH5CGQ5g2NtFF0gwz22/Vyqec
DDjhewYjm14Kk7ppiiWn4SYzbPHHbjYdEXo6GURzhZF5vF+qRrPXpoB0Igq2IpYcI33Dy9KnmWZq
YUYbnEt9UvBhH+hy0WS7VySjofOWcFxBejPc+8ddKPgjuTceXWON7YrL9nqJ1JIr+lSRhsFQw1LJ
6EFJKiymY9ehJ/U6jjDrw38nnJ8ZkTis0M7VMtokYl4DTukiiDpqtGYYNM4Yh7SbnhHOnofkQRid
2sRAuVk3tUDmE63Xhssb6O42qOHup3ohSNwZhhcLHnujS1Vkw04lo7gL8eabm7OoV/XS40iFeTsn
K7rHm1pO1Z5jOHicJSm852OoNJ6w1z3HBw1BKkucRPlIFXR5GcQIrQl08BSB43KDHammO+unihUb
31z9EhISHDGLNzNjyfEam0NvrlOUAoajmJyFXF+t+rVbv+4J+I0BWMUnFNR8btqL3/RzeQ8IYdav
g6r7aqAdbVugxI6SzbDXG+XtPRIii3GRjeQASQTjWVJlgFBntDZwljHSOJk3LtuJsLq2yhQXPSiu
PVIV1bxSgUjJBmRQiQ8XhCJ+W8LNLHkIahBOnAGabGtXqBl7ZyoLVmIs+LtZtW4uWu9UDO2ScNLj
zhRBnG9xiTFU5l2DgHlr2/Qm7xveVB4A/gf4djqTucFoq/m6Jx+Uyl85yaZ1GdohZ0vvt0xwfjp4
yoeaYEdncMvkN33+f9wnN2pkfESZSDGMzeyj4ZvIwmXayjHOCEPvPvoTkFCV3vEz3STW3su2qOBI
x2rs0+O3Ef+n4LtC0CEQrMQGUqSQsIZLdq00ZMrtSlapapZHxri/GHN69vAS62BPoIuJKYC+OFlo
Bubi17GC4YXQDST0ctlhFjkTfhsvJS26AFvmIZLgEZr2aIifWu7owCJA7IV0ibsH803JIhlS+/gM
iexxft2ykio0jxknmB3IZ/JS2RouyIz9DllLwZEcHR7iLKs+R4sRbYoVRBSgH4Gu2z06WpAyHbKH
9NprJK70MaIOHdexqAFdd9E6BF2CMOadMN1wi+C3chz2BNGEqVW0wufAfXnDU+AepkpkU2vkn1HV
I6zSiktVG1teqPzk8p7Bk9afI22sgd3qAzfEMoFCP5trOKOGj+j0SQRal9v2VIcD4rQnAdcazoV3
4KGFLMzk0yN20xjlaDWrQ2EWQIAvLEN2NKrhcr/jSuWCWpmWiczdcwrnbviR4Y7mpTy047yZ24/z
G/i82SzRf1MuojnxIvrJsXapd+Wny8InC6+L/FjEExiZgvmWH+JSNNYQ6NyL3jIAk567TJtS/7RK
BZuoT55PhsGaZ9luSHSTsRcpmy7ryHshz7Kex9i7mTi6VXh/hxL4D1i2IqG4exEldzB/CdY7XU+1
13XqSNNPqQkrtckNLPrtnKHGta4Tve3CtKser2AtjAwjIl6pLvqROAPsAj687LyaGCpAG2Dsacyz
sLxL+h430DAGjUuGx8iA9NBCwN05wXyzNaV66obEdOVF1IwTZXulK1xvUYWq4ZAv6NPZl2edBqQO
6B7OiXXSVR/nwIGnkTfPtU6felvQ4LXi+bbeyvgmJ3sG1Id5TxTETph5Qleaup/CFvv66yORd+xU
XIhXy9nYju9jWzS5qlmPd53r0LpnxqujIBrZAfOqy3AHe/0+6OuHWqBZ18rvve5tR3C/3ZVpcYkD
WqEfslj4a2Q+ZEepykSA+Jcf+URg48fea2W/PZ/frWEgpbmOYiHfW3qOXZ/MIw0Rtq2bRHP1KEB+
4E4BLmq/CBP+p3Ppy7jFS3xM9zXhja3qYQ/FrVZRi6Z7GlsxafpDIeHPSoUSxIeo6lVHKfRQyWJw
3LOLc+kdqnX37GV5K3M8rNHb0YDiRaMe45v7tPSLNkhbAKyZdjyeBs2THx0EJZoxD2mLOYsnbXnr
cky8tRmNbpCkBMgw6WH9cohZOAorZkFVkkL3/kCy/LJmxlq5B/hDPVYEQk94NCk5sK5QxS+xDUCp
iAPtBRv+N9exxPNhRueB68VIkE6H6kMPdNm38na/7mxKzYX2Mcgd1/PCkW/tKluZCAc4Zc1oCytZ
jpNVCXSfAhNrm1q/aDCIs4lb20NRgKbNoid/6UgNUx6VOOhFZX0x2ZseH0abAPEarsO88s3aHU/5
6/fqgj27BaAzlPK1XBGZL3+Y1JaY+oMjTL590JFanx1hQsVfkDz4EVtxQHEVoINBtm5+iVqQ6ZPI
QBXhL8JvWDRQDwchbABTXJmdHlVq9TVUohLsK0OTQ4Hsj2kTCoO25SwWzZNB/sicrDriwN7IytbJ
Qilzu4EFlspP8RiCDwBNmXnuwFMHuB9d4oX0avN4m6sXXLvDwExU0aFABePdDjXwl3GQlY4Fm2Ho
sZxHtcpyWpHkqsjwLqwqeN1lh+hxbdJA3cMf+O/OwseILIkE+8Ff4OvWYRZacAxGvafVcEU+z/BX
dEugzlmcyuKXLwzNTvB92cFL3WjFhcHRHI6M4Loz7fxXSHL4JR4mKLgP65TrpoNOa7pIxVIhB9SO
frI1DtToDCjj0iKnXadsxhYISy4k5BLTFqgVxbQyj83YD6E2ScDkWAAbbTl3LiFnEZZ9QgxbpLyD
c3EU6yzc0uUisfTletHE5/XaG0J9Tpdic+pSnacKmATs/YthT1qGUvb5FnLM3v9mdEXdUH/PjkC1
1bc5tBTS0IHrZ6ZUE5dJfCHuJNEdd9TfHyMPPSzrFbxEq/kH4DGFd2XYTZqnAjefU5R7MsjkWvQ3
5e5NviGhaZrY1aW3LTTiWUnyH2L96x2vyqheYFQllcGtm3GVgH24nNIa2oruNRmxZg52erb7TbTq
GHNgTz5Cm4GKgB7neXgWz0+UyNlTJTpaeXsi8Grs+qbjIvOJA9RwaB9ldDOAv6Zs95gNqPDw3pSw
gkQW5FrxObb3whSyPgKHaXPhxCuZNfWSUmT5i7rkuTCtvvngiluY5NARiTULFFnnvhA0CIDEeuQB
iGRoe/egChsaZ2bG26Ddf/XyUpEjD+t1ySWWAGTesqjUj2ddGU6IKTg9Yi+xyLvJ/PRAd73VvbJ3
VNgbSutZyBQPUQkHsTpN/Rfdu3mwAeDJ90GTsGqzTYw0CPMOCF9l4LRruwF+4Rh4MlYJfmgPkRqg
PGmuZq8zJhPKKm+cdZ58DZvfeWX5qZW0MShorHXm7NJQ/UnesyfDVSifDW7FXiPmo2Jt0/XYdvqo
gzcB45TPaghcAewDNtwKQXiErjIH1IPTYtRoLpon8IJvmMEmLGk1RPB5zxVRTBP8LKkpn+IIh6VV
4RCST5yFJsufLsQ643ZNeHfBvP9IitZnDOtrM6FE8rLnm3wmkF9G4/x/fFy3H8gmQz0RdEo2Eg8A
Sz/luHRe9DwLKVG+kh1HRF5uK+oHDeYcPebm4J2g7pxi/FmDhxg2pft+6vBCiB3emEgvb7A5Sk49
OSJYw6In6vrh/l509pONvLNm/pzEEifOJgkOYsQMlDNXMT3sQBVx4kV/cOUpbEQCrO4F5gm5fJ3k
ElXniyod5aqNP19BkOCUDMQlj6Byh0DYPiQIOEqswjKQCje8duQ2ygti8REcWUKEiy3bKfKxTfmI
2TC58x3Q4y9VIzlZ/JPt1TwQtEF7bYRRVyVB3LeKEijM67yZ5XClUG/mDPtk8zIDKCjK3b8uGXqI
OjouspQliRM8RRE4yqu485Owh6mDDigX1QRwaat/WFFtHg3/UDeNuHgRIr7yzgqGSt4FK6ukeydK
kdUu+FI3NHGsF2Phox7tzrDxTYQJ2LM842Q0qqEAqaWOkSlBvQ7eUaVYQyfR5mTAJ80RTrmHgfig
iAOBUYpuGvDRNET64FAGwJbzcQcOsdm9fxIBYjrXcWp4kmOif8zmvOU1hqFaSnKCFwIUhSp8d+Rv
M4mPV4oyIVHW0O2NlKRDEBawGhsA0J2A5BeODaQx7wGafg3f+SwtZYRKzZjPdZXRdP5Qm36yEFCe
I7SMKjiDJq3PHraNPQDqhtFW/OogyqAViGBPPoC/NyeM0a6ZKRdbvr2GCmbOzRMjLF9nZ5kDPeLc
IbhU6NNDIAvJmVSQ8DyPYfGFOq+1N+Kx3x+S6+NWW0XGocKx16FwlbBHbigRC6XPTDTAf3hH6aOR
HoHRNKliNHM7BaaUwQnRUl9veK0R2YtREicoUBoB/s8bViGanPiEk2rLEMWPfF5z7aDlj9bAhWwA
69n7OIuMN7StKmzSk7ijWGqB9GO9prmdH3Vcrud5RhS3TOzsfdnE445wQOS/l+EbBUr68kLN2jXm
r1jFEUAZJxxRWmV6zmoak9h9V5FYFMDLCQR1TZmcsSjTlBCsBYGFDR7+Xv//ZvAo5EVTn4+ocvG2
TSHDYVTIFHXds212k09mv3wUnlbjHFXL4E2btFuZ0jMlIEKHe+/B94vPy94LCThduoii8dWaHopK
Zn1OWEOPwR896OPGwYnHddNj9jrsv+Ib/y51V90sSZKd8M0s5MFHr3SLwjyXG4v3diahdAv4f6br
u0ijVahUZRihFEKEZgiHpDN2tupAmQ03Sr0ljU19AZbM1hNGrqm2oH4eih0hTufNuZDYHr3H4fjs
HZhgdKWyY9eKAYV2+Y0/4Wh/nmqHrfCZ4JwK8OEDku39NfzePDKKRtGodval/7b1wp8w1Yty8kR0
DSICbfOzDk12T/cgQHO3yu1mBlEvNJcq+Pphf/6U/wPh72NEqhTh87DJEqrPpWb0DAtI081tx0IE
Kt7nY/QrLJDVIN/1pdui9WvJ90q97B+MlsEswkC3SyYLLEGmN1YnQoExsJ44PvC/MA8u1AUfP73F
UHGokGVADbQktuzQ0GlLIB5PbOv4w6qo1w3yJPNS2KY22HuiwkZb3sMHXYxTBit27L2LNI8FvS+4
wpr00DR7iR7jKAgXEmIqpNOtgnd4yt4EModfTaHK+xqZwVNrk1AON6Tg8sziOyXpvDB2WCTSOkgV
+MV0caR9zB0ADj2ps+4wKHEqQwkBB8HYTLVfup8iT2bqiaWnThH7qYDtxkWPZzGSBqAME8I07Z/8
pBLcGaGpxGqLOSSY80LTk4hAFScheVegM4Qm+P1UOi0yr+jWm3keVDTQtwvhy6Uu3SuczNWK1ieP
DaNF4zlXI7YmttJG7UlpVpV4JWzylfc8LIzWQnEnUDT9pXhX2oGMM4upYm3p/wdc8v2VeCyObikz
iCKhcMmOEdrLZCfwDeZi8Vjwz3vEFFXTcadqd/k/sYQJnENNbDXTgoHyWAmlD4XE6qFTJu6DpVKK
QtE+DWkNsZGGOpPtDxfUM6tx4EzF8Qg97jCredgHYCujua5DV5hhZbrIjC/Op2IEQ4mfg75rsLBh
pH87HzDWYDdpI1MObMe8oST9sM3VGzOQItRbnCDqaFHXvWhSxz42fjeKQyQ11bMgNSMLFGFfp97p
oTLBKXeDu33k9nXguCa3iZ+FPDPaH42bsofDeCDAF1r3LgZgjER9hP2Pxt98pezADLI5w/N+eo7O
O2N7qjxnDHUtiwORTKdhpcklC0h491SNii8uCAUq7dvJ8gDmc0vPq1YB/LgiDX0FGs9uDtw4fv/o
mPetFMWWygSp9A3hYPUpmRAkGJyIW2mLyQHz4bB5pChhYVx0cEOZ/l676PGDP6Z3/1u07/VwM64M
ZucEimpBh3XVaEERdml5gnkL7zGimFHXQU0yhYb/qVlt+pkXOISgS6Jpbr5s3sn/3295M5sQpg3w
8kN/Y5Hj2yHpJq8ihG/JTb38yqPz7/gNqlBGklxqwoTMasaoIwEdnVyt9TXg85MwpD/BcYpcNmJz
2mpAZRoQUDOQkiDupKZw19WvEx9S41v6Jw2hJ0P3r/fmGbbuVfcXvrlCu1xKSjf6u+i9vgzcOrNv
lI5uC6mnXbmArJlMG1rOR3M7fC9jhoOsalNV6cLJbE0IziUxMFZD2NLwhz/opwgK1/xQ4EW6QEa6
FuEPwfJey4GuR8rar0wR9249PkY7P78jm4rG4qXsHhcosX/r6NZXZQ2dAjY3uAPKBIatfWBS7z/S
R+LpDRxkrvRhY7TUtd7e2n0x8WMLKia1PyQPwATiuLll6DZ7ZpXqorvMRtPrU2UhsTdr6S1ku6iJ
ZG4yVZjWwH1OA0UgMnymWdcFOvpCjoOn2QlVW/9/kEJgT9FAPO7BBz0jXmOg5G7PmnbBe9yguObY
Cs542okjEk8j/332D9mfzKZtIprmIwpeoyDZ78KlFxyvpzcd7oNMtVUuttFkQBV2oRN2+HfHsSgw
SFsLRStZ1gwEEDsiLtL2y5fELYHNB2fDa59qEpZ9pytQIP8c5yHTxDdnak+FsMZqtbtF/PeUz5Ag
/1R+qSPEw85fwkJjeSYiqICWLHBQTELz5oRiLsO767n1tBsIaC0Xd7LF2ovEUocgMyCAU7W//jY/
BhevOJZ8bvdMSAy4RpRLHSh7ACLBK6MEP7Qq8VZII/OgA8kA78SfBdpa4Fs+pB3NfK/5WcaYAf3d
FNEBpo3wYtzpc/u4Ze241gpxWb49XsUFE6uw/oNTyGBCP6j6f+E1Pls6KBVvcDHGtVmkx+J6GbPw
0hgAxNTs64VhzgjxItI8NY+YKD963gTMP5JV1ejv9rz66XVE01lG4mA8PZ/kBK4i29rSox0q9nWj
X6Dq1OXUceA1XO9/tloIGDngV+qVOK1QOqix9oSKyHmgnpbzZ9YtapjPwp52NPe3kHiSSK2Ool6U
5DirVA53y6gA+daifLjIPGtknoXA+cYnh7GVv4KGAbQBhMTT0FF9ZL2eoCgBqIzfrpvn4w1scbE8
xZlFYWujCgaGRayOpm2E59FUYt/JXIS8ttF1V0BeXqkwqPHvSPm8HfzM1kv8pNSliz8UZtTiWiQh
WCW8pH89rQh0Jt8AyW/UyHoMsG/mQuL7KeWfXs0nxBVV4FRmDfrhC/UdxepOahuITTUS0fByF5q0
ZIauWHkqFxQvcC6y1azOhzW4L9OEjrenqklqFah1EXReEGr0lC9HWAkFgnUf1jFJWlQJJoyk5h5f
GORmZ8Ted6/zNDdzM7SM/YENhSsuJD0QEYxsBM0noQk0CqXoSxuFQ6eAoOzJhJnZ3k4LnEcabEOF
IS2zkPU0qrxDsE8PexqmBWd5/tsTTzQFAp57yFT4lg6tw6uWexlqmDoi5fAkRS6CyucFccHfVrBM
ftO2U8pF4UHaVtjiopHD2sfm3iKEXbef8/Phm3Coa/F2O6HqUdwCDzBqtLWyBEc0LpLi9PWIHOB8
PKQ85BxYXipc1p+RFl+1cv4jQQZq4s9VGLheqCpiJDPsRWmaRTfMseEd9hmsjrnm6fJtv6KFNfZg
O949xrHPJ6ZRJpQKKBeybZ8j9RzwZJ563Z/oxGeuQbXyk6s4YI479iAAqHW01ThJ28xQiiSetOkZ
QxyncKXrtQiFZFPb8RE9sY0J5XALpjQ//k8YCikzfsahuj2e0n+EgVQyjyI+iBqhIdvgF1XhcEkM
O+Jj/JAJHomMw+yQ2zrUovkBKwaK/4/WTAgEsJUpd8QKiI38xuSWxHsBjbroB9QDFue1JXzP3h07
aXAAoIPawNRi5WrEiErdV9J3+pGJYNF1T4BdV8gdVhBejE0mZRaHSBiplbfLqjBb9FQuUp4Jm92X
qsajLhl6Migl9O05/ck5Zgw8kIIhWK2EiG+mDKAU3rIbIXtiRAc+3WVwierEkhASIJuZ1PGXAS7O
6IEgqkypUMLUE7FyJejoLyzZquIGsH0tslakytfqV7yeXxeQkx87hDZgWIp3DRfGrydoc5fILCzp
ai9EMnl5YoGozRHyLRlC70Q5YEds9peqR4k6O3ob+/zaRrieYZFhl/VcPDCdLkXyuE7gF2OTMEwy
zSVrC1SI9N4u+4AR/D1n9DM3Q/1oAnFOKzw9D/A3kdNHxHmca1DfD3uX6as3I+mKCaeNvnW8OnrY
3XfLcQjVZdJHlTtmm8R9D/Zc6tjRE6ljlluGLkrNTgJCmhjfrpHtR8LBnkQEn5m1yDpj6G4iZFWX
Q/8p5Y9fkLGTnjPyzJtVrLUXFjku0h+/aFBjBKPc37JVRmOXO9BsubuOXvBdVt8ODwYozCs8ZCjK
Pg73UiX4bLSg3K+tgQBJXYEYKtFPsS/6lKPjTnOwINM0C44gdnnB0ucwdgT7pXy0g0qvcpWceDbI
gcor82q/5LfovIW7Ve/Rvw6Wxz2JgEjcaSbhGtRVVsf3qIZez2gqx8bcXmfpUGcBybtSNL4QHJ/T
pfh/hEEpIz9pGWBie0XQeEoxHnl/NjV2Wm41wH0T2yoCn/MUZ0uxfht0Dkflf5DZtJ6aehniyk9k
ZlWqucwEgsPK2uBlI9D1M9U94tzoOp36gdqY1KQCe0JU/Fd/w+D50GjtQJ6VpLwVm724qeqS7M8M
fBuuDtsIyo452YdkCcDVipc5VQhfhVrFspmBYBxC/j0a3BQL290Qtg/N4Yebch58LXkz1927Q2sM
Mwj07o8O8kJX1/7Trmc/t3PKPh5gXO+fSj9sMGQGTCJ7nSHiBioTieVEFaG/gFL7WjFC7Q+1806B
tk9slXiXywzT4aS7lDImPkxBdFRvIptY5S1VTMosGLZiHJNgNRvDgVJ/O/EtX1STZnfvsvGN5D5G
M2dYKuU5cXQ5IKzZEgdvUC1iHEH5jpw902/Xa9DxRWlXF2T2+oeHJv0Vo2O16a+On44rsRP/fNXz
vlJNbvtCDTb5lLimrq+Z37mEJDk7202fIOufB+JWynWutfufSmLuuD+ve3jFKEcsbR5VIBI8y35R
o+s6LKTJXcHdOilE7wMkv/6OJg9r6aJaMZnJuKaLoWZRUog5lq6SGClhgg0Swms8UlYY1Sh8lvSS
stEuUnRXdEWKRyHsDvMel9m8kOAR2tNdNGMVHGGKHLdp+B9oe9EnnnUF2rGLH8V7K37k//pyE9LO
sQD5lj+2BUYZqS0jKdiU1znyMyqirGN4+s3rz5/o5eGXJeYVAaYhuFC94e5GO+ChmfIX0GSWTuQr
xFKKVIyOBz0gMWSPJ3vlmwLeOScdXVUbYNpWvbglfyl3xoWkwa6mNzhovZVlBwZlCkpT2mQxChls
8qrL1HAlAE2CU8e+CACtxcDaeskm3pKIY9UHS57EOmJvGEcONp0xY/73jvJ58U1d4tW4aDuLttXr
wPU8UAvk8B/Q9QqHaFbmZQxeTYcJF/tylLLnBcjkUeWK0a6qTAOMsddx0Oj9Se4EJ5ALbE7uJrRs
6gJVLq89xGN3KbsO0AYj9/fPkHJ0yWaXVvrsDl/HQwicDzMMhGHSh6YyDOvwnQtfGz1gcBNF/HtU
EhevaNXA/BkNxi7BU+vMAah+/ACsqbxM60+PKCcE5Won0PbuNYKPuhkn4dyUz8ce8oi8Ykdc1LEX
9b7ZUrfnDUfBJ6aw73DGnN/6P5BM65qw+lDz55aXaWAYPrOZZ/N5ZeLbeB2w3u04pP7GxXbLamxB
waiW1s3unRdiQBOurSyLZUZuX+k63la/ItOG0LWRNHwxndKgxuPyvFR/OLuieXUjMI0Zt4cVInmD
cJ3lV3bQyOlX5Ru/qi4GFDU5gBWh4blHLvX3c4/sOi6xEuvVTSouALVe0uGt+8LMZWIiG4MGRfQl
alu0fdKF6xU2HDGfgME48dZxo1l0IW1vAHcHOvC30qBHmF8gkewI9wHae2Ynn4GF6oHFSMe/Ei0d
+qk0p7CqG5Jb1atrfDm2dOk+fl19lwGHdZKZpYEBdYtgfjmm3YKXVEPM5SkCfRhK+qPtR12lXDSp
knWPh/kO0FuO9wmeeQ/LDXIVbqsQVmv3+cdfR1JOAnQ85HERuOAxavBif1IZmG7sI/ILRl5z4q0a
4aP7SjOjvdn5/NNru+UbFMxM3AYNkThMegCY+Skgy8TjgsnEu35WvHZs2yBWiFvW7ft94LgvQWpj
yyuh/KZ+zO5T9216cYl7CeaUsqng/ssYnmitfRXig9gXUxQC3HeqAqwujbPD6V0Kz0/Kn1D23Ihn
mbd3AXuRSdnBTpPyFt6oflIre6IXYfqgf5Op4WradiDL8mds+9eivCCvJj1RYnHpwjZnl2ieKs8e
WIB0BO09OcsGNDrvL073F9ZAR9Y3KdZeWdm1xUtmO1zMdJu3IoGgmFH5EWLJ0b7CgEGXXMT3xBru
uywdxUluUtEVoord+Z26ygTbh9KkuYDqmQuOZKDCWcYM83+RKmioy+SGyvgJuMZrATm1rbAXyhLZ
GBM2z2LDunRGk59BUlSMGa62whV9Y+6ZRrw7xbbnFVRV1wFGPS6UenFfCA88vatcZ7OeFo4tvGQt
xcI/DHkhrgsOuiy7bfVyczgxXAE8tO+cU0yFQLyQfK1LYS/dJw7MZVhLzzfyMXznVw5a7ApTgB+p
8GMLhJUnxJeM/sqrHK82YZCJRmtkLTdVoCaUvovzDwEoxio0oHrAxym/lH7ES/Q79UHZt7kO3cgA
+SxacRHwZKEf97OyTFBxW1JJ/n3MuAauXezeeiQhVXswItae6542ycTchBlbVN7kl7rSl9sY4OMM
InFo7mKsTpbtZso5Fr9Usc42d4Xro8q9ub2/1i27tdIRJEVW8tVGXpbS3GsxKBeg7h4QZ9YRNnOG
nCq/TWjTNEHTSsEND2k5aolM3/yMvYbri7dkvadWRNLYMgbHiRsgHBx3m6UqYt7YhfNW6kQnizAo
9AHLZa0j0/Cqk7RNrvMWQRNGEtqUdLHiy8b8IWgHNmevXU+vSH9HeC+/79Ut8zv0qKKXZa/UWEsn
nH+4YbsfTi2um2sKvfL77kcXF4/7V+0kOtuH4JIlpeM0Sf4HDlgl1cuzkfEPQISuvucNLcAyJZE9
5xI+7awC0a7qjDG6+5ja6BEbyACUOs7we8bNn6gLAL6zC0bEXdX6xb9k5Sd/7CpXZ3T3yroN7EIU
XPt4WoGCMpnU1PyoOj+oJl4RipdJPBpxSwz1lD5zBda52sqwvQIsBkLsRsbGKeMJXcldF5K/9Wbh
O8FgX4955k7ze12jGkqfYzRHchbgOuTnHrsbCmB+4O1ydWNTuekpIUnq7JdooQsDiiODBvAUnvUB
5Ar+4Y4vsGqkZepXor78zn583oRs5IEP2ja8Su/qjDUspVCuekcfpeCQnKLsI8GwLU7HZ5P+1Rv6
vGR2AL+ggP61+WpJPn/3JmFFsn3BI/LiBDmU01m8nZlu/Zny3TkoX6obEBDV27dhr4KNNoJW2Ab6
/hKyHQTE86XEKMQOZxn/AmuUVcvve9PDDkeBsiaweYwVXgNEpxuHGL8IwDpXI+QAC5s4yQz7KNY0
Uchvr7n65n9BBL4G17BmAnb+4HibEo+mZRZUYYtdtaRvXZPcLYLD95jiB6WLkk3TuELsiOFBi8JC
jsOhpllAGu6mxMcz+S8qMXm0ShYdvKk571evy8Uzk56RPOL73l6HUfLHRQ0jxhnxSMQ0b/c09M93
Lv+QxwxRBSrwgZ+ayT44k/exPnBAAhY+KzIUYRf4rai2uQE4ay05HcLpPdDHPaCO08lhvpVm4RPX
KYs196nITdok3hPTWfvsCotku26pRDHYWhMbiCzYtJyL35oKBdZPJbMFQ/28jec8sJBH4KVpn8xj
9gIyPQsi0Rhpglr2bgwaFgm+fxIfm1K1d+6o7yMFQOaSb+K2aSTsR0OxNPmCfXmbey0+/0gyZYU2
2TGc9TQCNzqxBmK8O3CGscwddjiCqBLePvz9sJUx2mkOoCJtCAYv1UhHWRZbuSzkuZk6i108hBff
r7ixdKkkhUEGpH6MoBDW+D1B66e7mvvUENL/X26hzhto8bST4GXAgcGQGGBm5qquuUoUfEs5g69O
Ws0QaPd0DX/emRvwHB5Z0R92okpP3W3Vqb+3mJiCBon1tcCj7Ry2zrG63HAAIpYpkoYDkPUub7o8
/wImSowDP8EXlvZJYK/J2RURtoO3EvOmlT6odFZ/mg/5aeK/gftuE8XxCyVc42O6efD/mqyoWnC4
6Wf2M8UdN7A0Wcq2bFP0E+h99eFQkiBpW/Wu+wT/JJSaKu5MvZl8A9cg5n9P0qi0PQ2Ss6/KldNQ
KQn4IsYTiv4mWF5tzmRPwOUv5Uh/40BWjGfB5NqNFwThLFHAfnpatw0PsWD/fnL2/54OgC7QA+EY
ll8Qw0x0n/EAovQVIdPfz/rGHbsbkRe3v+IPBsApdPBxA+HTVIC7cBQkvzKMiWvV2JxPejQ8a9o7
J6Zs1uJFl+m7AQJ1SX0LpxitnUF75//VEuTCW2X9a/WnzAVLnplhY6h4euxi3JRo1W645P2EGKg2
slR4GyGwTs9P7t1EYGKZQuydk0k5tsquCu6vFNwdeHt+CuPupRy6XCPjkBZ57h4pbFVBNSseq4rV
zGSe1rT7m/K5Luh0hTcbYK13PPlgd/FCCnrijA4tRDeBuZ/uS0bIvi0MOD5MrM4DOeykdcZ/79fV
HtvMHGATIATMpzqrw9wWF5EpsliD7KKDlM8KQiUhwItq+KrVkM4lVfUgnK+TmGmxmo5Xd6oYU7MZ
huksFLk7uIeuKc+biE/vNLJYDtfBv9E/jUSGjXYy9Lqlt1UG3br2I0oehVHJnBwvgugrymR+q2sa
Z8bj6vRy2jMAjS019levtkY82AjleuU0kAVXjKoIl5UAEnaFYYXQh/4Qp7OKOTpVfv6MqJ/Xe/8p
0J5f3Z1jnPbRpgpFLnz71y230CyeXzOjl2XpilbWPga3uY2iMxUOCj6ICNcFgl2pyAsuS8UCmN0d
FzZUw6Dzi7Me6to9CcmwecSV+UuHWu1BG1b/PCIThug63qIBo89aBREfYJAtg32JO5e0x1iblv1R
fmVQSzAqmrMVYP5qKVIu4xwa9Dnk9zoRHEnyYSmvEH1+N1WF7pJPRQa3QSoyA0REv/vBcPdksTO5
NM2CtzVhf0tWv4kw+vs2zAuGXF6oI2CXjOa4C6I/3o5NEdITh63D63zdKTOeKQlPVq7o2E95RaN7
HcYSjtkntsddf7EICJnzju7aVDKY9khfn21KwkHBL88Fb7HKWRmdTgepeEUj+FOW+PzqwwGS7t1R
BppW+hDMjvjJmtp2qKEVObHtfY2XIZbY6pbrE5VbK7bcNZ6S16MaTmUwMg8t4XCGeAwCvbNVnj3k
xWXOZ3GINp2jBMRJ8uUzG8CcInJH/cyrKwKtNpndaHVs8COcsqq2CQpDmZ+Ppq72HwcuHqEwuJmr
NodmLudnlQG41WgP8dIYrvlwz1kqjcx1e8Cq6/gIiEK2xVkkU7AaICJxzypbFEM6KR4NyNjVchvU
QbCan9YwWr6OKnsTzW23TeozlxGvDUGOlxovEFWvwCDrJmbAlqt01ERF0PbuTK539R4ZXj1/U0ei
aURaaj2UI5FtZPd6+PLOpEX8bYby+M5Gosma7cpmq0Viq1XEdFEvkZBt7lDzxBjyFYL7JKsWc/NB
n8F3DresncoIxWWfCGtQgR/kNfGSStdi5Xft2/sM9T45lfZwV1BdPjmuGuQkbb0IEYIbEra9msw1
I9rXd5ZGgn6CbDwkdzrd++Dv6sTpIXni/9tOc1j71snS9t6gT6hxZwOrvtYo/BCoxH87KAcchdD2
5+oy/Idm0jG8O53GWYEV6km7VWHnc/QWHSJo+X84jqxlIllUkW49RB0Csnx+XTgxFir4PIMguTtd
wg+HuCkaozDldq9KsUVw0giMZxOSlBm1QuutGkra6R+xcDagDsC3dThdD9nWv1LBGqERMJRUFTxZ
A0D3VkugjBN0G445DUAobIhhcSscj2E3iL9P3HW1u5vXsdZj2tyzuo8R6fZvJnJLkm7J9yK6I+Il
zEvUFhc7W7cO0oTmvUL07IRb47GL1YlAkcHut+dmaFY99Pw5OgycONEE6I0IeMF9Q8qJSS2hiLHm
WmDtuictlJe8ej7hrySHjEIIQ0Bhs+AgO2Kqe3I++PH/GJPmq3VUeueKhPR5DaeCtvyPen2fOL9V
aT0bhnW0stzMDdRneNXCkDN9iDZ+S1BFpiru1vfVK1ud/eo7iawU+1KmCi6mFW/EUJ/j4SiDlURe
j2UYQCU1mKNZ/L/fMvWVh3PElrpyh6FHVb1DPR40heZPug1wlubkZXwg+ot+2Kc7B+3YhJc6mNkq
4q71GrQoUzF+JF59NyvWWWvDk1QfwP+xB0tmZy/0LGudArhLdo2xkNydsX+tlf0DAflJD7GPF6e0
U1GwOcGDwTgMjf4oC64YbRtbG6lVNVsWi2vMwjZE5ojZQrOJ6ACG57EhEcXKtpd9xJ6x25y0tXiv
RvNiyMVsyVSv09fIPt3jxpBaBhILhpsIbrGZoW6xWY+PXFal6yCAmJiMx7/lyjWhFf9eK4a2WT8z
NhYgmcaml0uPY5owuINovzwiVOnDtjN6Wwl/y0IbXnc3i9Z3pxVyAFqb+VC7IBM0eGfj7RjplxJ9
GiKSwTaxPMJUzYCl9NsFiNfSx1x4wqILRGeMzgRNoTEmtBT91MLUMEfWlAlrQzLDBN0r6C8HDZzr
k+l7fv3AMylcIRG/VofxoUSTC5fnZ/Vo0hJqX57MezmL43FsMWrAYImie4xXNw4/YOpxw6QudV7C
k4n+1/+5IthFgJt33/V+Sysl3Vv9ozWzXCsZ6kddMtq6CJUESqy+EOSEDjtw7F7nN0Skx3Ftq1dG
rYaYN5YHsxUILLYO7DJrla1sJbYzmEs9+KR/CyUO1EVmp5AIdmNqk6QVkaXAfdhlnlg10wAQFBHE
rqZy6Y5Fltsuc/TaPZKca9NQFtHouifwjGyAb40MB53es99mRAAa8waJhn7J4v50oWpTJkrPbAde
dUkNjQVKzUr6NeXh0kGmw2uQNf8+R2uPro1Nfi5tvjaIK1q48lllatdPBun+D66kgqjeubscfrhd
KlF2xvOxoUHiAiWBEHD/RkDM6DoHN5KoaiuQmzPK8fsz+cyJidoXyPKwabxNAX8M8MlzLSwkcJll
esGitnuXtlw26YSZ9EwXq3QhJ19MdFc6vHfSSEJM6zMB+qc2gANy892dRD+SEzO2tv5UzOIqLVjd
wbS+UDB2p1lUvqmQTb5oYpVMqHvxMnNm5epVhT5J3ujM4t3OZcCC4+2iZN6qAQB6IUaqeI7rRyNU
j4LUb8LucI8KNVIxk8bzGII+RvW6mSkKXpIj8EGLFTNSwPYgyn3rAv4CWRHEbBCrBBUWuf1qJZZE
l5sud5v7ZHwMRMCYMvzz9WGbfMtAK4L5KfL1sX9ThwanXQmNy1ivR6PN/jO+3Rct1zAUWmodBYsg
DV3UkHiQ+bDxDRMhELj2iqYfUoecfk4Bpq3wJVI+7BBqM6eUG+qO4aFguBYOIHEF721Ws2sljGlg
RnzmvsnR03xAcnMX74SP5FGEgIVvEtIaOwdBk/0kaQZ8nfiEbDJ/smzKDkXcb1Y5sP8uPh0MyoTe
LR/wgHy5n/rqLO0B5Kl7XkN8UI41bHT+lz4U8yZ50rIsppw1YeaPcOpTqfWh1f+vFXUjROdcwvGc
BaU671WJ9mga2P4ckbv4qUiRUwuPd2LW7ncOPdd7erBAM0Ll/XoE8bdSahsjk7Z1ap/3nPD9D24O
7o/utUvlhoIM5WCTGLJ5Dkq1M7ZLXLP414IyCEV25Fd1qdQk4JNe8NkIf1epVlDiNJLMB+oisS1S
qk4gwRuTzw3NOJKa5Hxenf9fhpeCjhBxJnqVHzaLnt0GCKiXhHmiLK37G+AvzQVKFyCXZtF7Gidy
e/Kt/YV7EbtqMrCt/pVycLZJphCw1jn9bAH8zBR8uNka7MDHDFpT8nsQQTDJAXSpFWDN45b1qceH
TI5JpA91E5q6zqzak1F/vSqrcr8V/OU9zMSbLX+JYOqUYie+WE0jKWKX8VnB8W3sU6Wk8rA5JZ+N
TvczLqBZQRSOn9gnHgDmljx8Iq7uJXidl+itSahlCCzZXzEX+jeO+PRKnVagXZdmOcbXrI25Bwcv
f1tN3qKguA6WRnaXhROqgdhwUJtbm+pwW/MUoSqP5vTIend1JrxMO4reSxzSE9vHABjo1BKvilby
RU9UfFLe4+Gnxdn9PzMWg2LUPPNLSOLQqzdDis0QIY6rGes3chAnKRkclbSPrlZOT7EH2/PnksuX
Kc2cC5bMPnp0DzvAX4pTwkkIkGdm8mer9L+x2nWj39pXA9QwpLNQfc4I8FiZ2mvNerXBFia89PNt
iNZ0Hz9ob+xC+iwH+2gjnlFoNkqQOYd0Y/iQrHS2OkBcjhsPp3ygejR0KoiJBPem/CQM23W+Qq/n
R1mpsTegtY29fgZb8y9q85SX+viD3gTluTMU4WcQ/j4Au38RajQOuv2WW4bjduXs+APpfHo3gvlX
+noD3tOaypKSrZpD6JkVA803kuWY9/5EDiZ7CtLlPfeoyNeGUQM2Z79Sw1A8Owrpk0fCc2dUGFxz
reTh/MTREMX0pL5jJUF3u4HCa1VPWiaGxJHGmgr58xIHVmxRXIUj2KmvvYUDE7BAxY/uWgkBjNVq
H7wmJbkWeLIgVJFBcFXEsZ/oJqwQh90eX01ja9SJKFy/Qa1U+UJELAzSZBy0hkmMbDbjvs80QPyV
hMPtOSwQdrHvePjqUptd/I96abv2tAJfulHwmSKW2ueXM/Bg9Kqyw5T+UMR5XNev4wmVOJcQoiXj
Pb0J6CPX2lt9rRg+lIuR7X9mdXCE3b9NtKPpoxx6gp1xYpzg//NMa19zdwhK5Ad1nCuCWRhkP4e9
dIYuU7d0P1dPH80sfDM9AVc9Za1Te0VOyO2RsSvYRIaFb7ZKoX4PgfQgKsuEmq/cJkk/eE41CSsa
7tCmXscjklRObdAJkM6Y8C2RwmACXDT6XD5oOVfsxVMphoA6V2kT7/hYxd3sFLRd5/zxyALf/j+A
6PGBkEq48horjwRAHbfZheelZINMUM4b5QetqfdOhLKeFVREr3akWlE22om3aDSjAQVJY3SQGhfm
6m4Rl9ycTGB5EycbVGsmbj4XmIvEQxa8Cr/Z10m42U/G0I+3BDpUE4X8Vh10faZZmpXPgxR+TBDv
o40h82obDHn1bzNt0ecgkcUphilL45LgMAunZr6xQKgGAN9ARPGbFfaQNR+idKx19YCUG4TE9xdK
l+6OpLGQHa5L4kw17BpsUMxxaaw0jouchAlK46GONipC47Mz3wLTLbgIGqFJxM1M+pRYkeGUBv20
+S51RO0r7eLyN/IJtOmNC6qPgB5GQ9mmyr87elWZ+o664hLaSdCx3l66UiqvemZhylilhBIzXIbU
i6WkQOAig4XnU3hmv99vxBkGLM1+v3ojB1r8SZino2vt9E8sfS+65zp+7K2jB11ROzGSrQBEC9MJ
kC4gmBVvkXZJ3YDINyNdoZrHExcwRnkDHoXBH0da8RYB4/yl8au5GmmQjJvRCMvUENmiUTbggGUG
sqp6Xkklt7QgTqMH3OgXSvrGcbEDAWDef2xYHKLjUVHGTx7jaFDVJHurbtKu8zctCuXORDCYydAT
9qN3W8gCjuGpj8izg2BckwUDo+dMoq+UWGYLxgqzBc4dej7lqQ2jFdgUTBJ4j5g6Vw5puGGDdDb0
xQgZAhbU9cxH47zxxIBy9DUNGs5YTCppNFE0ySpjcPeBLLcibCjnnH4Hy2S/QNVVbMzdGFOeFoRd
c9nKqakxOAXUzevdO+hhO1pfOXLOeOymh40yS8GTcv3uMS687pSTiLfZOUD3kQ8K05WrRzS708lN
nWmfTfKqDmCipYPqbYoY4m6Lu6JURqNLT7B1vjf+J6XYcuxIkbWPxaWGHqCFOAB3UTLxwCVu85AW
MFN4Ev9n/u6yU4z0l7kXRhQ7iqYCumSgrde/FrjXLGYm/sQvtYvMGyuNDM8ORLG41FgJBRf5+5HE
5Pzpoqkvo6wcGH/pqELsJ1SUrpuZ0/O5GHl3kLFiqKGTOTZsukP8XwSJ6smbjM6juv9vhRnB8VVw
/JSukir7NvgjCjag9dK0X3K0rfdipyw2AbpkC1eMiqwmN8z75wVRc9/H6nnkZG461BqE9gRJR8CF
e9bQ8VkugjwESh8/gaRGC5AvWrYQNiHuaYvDFj1mJKrO7cwB2f8yffFQHbKFTT6vdzf9bv1FGIdq
LvM6SqEmzejrP7xV7HO3tY+Or0cM0HhDVwahuQqBjbe+GydaDBO6QA6trVVCjd8CUNMhGzJ13X77
BWlkoSoynIF6WZJjHbVC2wAA+IBzhjoUjEPR5JOcVha9LmCoxmq21qpLc7STFrkeP/CQpJV8B8/0
McUsnEx75swnnMPmzeOQrb1JOOKvwrh0g+CCElWcSR1/VplNN3mExF9dEgpGmmQcV8pJYUe/1gEu
qSjexqGcxv3hbiEACwuRwNKjbvwVjzGuMNDg3gWZp+yOD6FqwNEhl+xMvtyP+LQyremMuzvH0zze
VToSaev8lzGrUiZNW1qvliSy1WhXxoWMt1t+x2z5LgzpgDd3EHLBuFohPeyVZDznMIoFPtps9BME
t/ojNN+oUvOmfrpc3Bfl+mJt/qaiWvxstpXomUIXSfPlQAYQLyaMfwvhiVViN0ZJPyVr9nImFxi9
s0Rz8LiNhmaHx6V2FtZlBnVvQR8dQsA2Sh7utP/QJhNxeP/ikcs127xZ6y7Tkzjz7//3nLgm2tYj
6ZlXG8Cvazvdy/AOJwieVQTPR9UNSuanheMY7+LMoLW495xfferxJQAY7nUUIc6ShDU3k9OPnqZ+
jmMZQWY43FDsUFKJPSKtmexZX9thupn38tKh9SfFrfQ0bhlM9BHUH6Vn1lNiB0OsToxXT4+6eDhg
WV6y7daaR4DjJk/KkxctQYUrbUI5GbdP6VMVq8x8Uy/UtU1ey6XaCOnNnkNKPmKoUMuVk4e0E86m
zmJQ6oSqgIk8MayhMQM07Lb0X83GWOtGdSXuILwbTzd/rkgyYwkuv+zG8hhvDeK9ZWK2M1cTED27
qZAmJRQoEkDQkmMvMrGXffyo7+97/TIakqX5un/KiWygtNiv64z1Tq5rESDw8t5Gg4KShk5Gm5/t
dqUTDun4Ag+4LjlC4piOJbCiaIQ7D91ofaJQrdj6jjIZ0Lk5CC2a8v4kckX6gSxNTC1jxnjivO92
KJTZ2AI0QFxuBSzzcotwe5o7in0caIwOOtCOvNf15jC+4WVUf3yQ8O2f032pzlO2M2uxk8L99n1/
B7e9XfhsbiaAlpexBeUIaI0hN8lJFfpOs2wCm6UUra2CiN3ieUOQ86IBZI2XCReRJzATsQD2sU73
QdNU5WUUsiwVNKPf0/vwCH6QRiSQ0jotItX8ZSqigsDosCez0wJ6n1C/4W+m9EZ0+SerFheF7+P8
vA723lna7DkL74GydmlS/v3/r/lGCNcLr29JXCyP02Fpl4PTnnMEMSulsUaB3tCcLjBwGIfF52OF
VbT2vfmXc2H8LINBpy3jLQRP1onQh6WbWV1aYxnPMBqRHd//72YjdeQ8PIHR+89GuWFv/oV0v1BC
C5epjonO10nkNhm9H/v6tJ1oBFnlW4HzcA5zqFkDKe3yhHnODApcv4ALRPd1IGo4RLUzmao9CTGC
xCr8Bhc76vWtA7oy411wWd3eEpx7Pab/ART0Lf2bgZ6HNuZRuR4NKWVq5XICz+MpDDKT7tRc2gaU
+ku6l6MPmNLr43Cfl+KmYyrW2HND+B2+9qsbAjVdIwNpovuk2JCdqwzDEtPgk5CD27M0JmKK/XLk
M2ckNF2rj67ZHKKR1CQo/ABPRC+QNuH6sQrK8Xuh5bidIzGSp+Wm9HVJ1DvUgvpVxjOx6NB9j0Cg
ZJwyHJEloR1229dpiEt6u1X8v6pKAsCc76I9D+wnqQrPIwgM92gCRoF4rjWS6SQjAh3HbLKvphit
loBaCtxNSsN7PZ9nBfBM1kiD6r7hztRl/Y9wJZcoxaqc5PYH2lHQBxczNwqAfBoyNxHrJQ2hEuRA
XxFfI5aCPJpcnQIEFR47RhOI6WGRxxRH5lPel/AWkJ4FYtMp9nX87Nv5uQbYn/oAiHTWO3ycPzh+
6IiD0DG0+kSwWrC1eqz78z3Vg9Iemb6PR5NwX+poU0K66lfiywnE/UPaPzFRE3j778kKihZ6dxaF
3xbiz1FgYUucLCc1mb5UlzlnUtRRguCI0dXASMphUUVv8tUInzO4QxAodJ16rDhbio1lxzrHLLNw
CBCaHA91bPwrF16C0JHD/bGXpZ4aqNl0ZpRXFEh8VyzdlzUUDvaLdWsCBLNkpOb/uJshNuNBs0K/
eZAXgjKNsiBoH/wEH1uKm1qu5cwUDc5kfP9WrmOppN/4BtQGRU1jp3lwLA17hqW7fmqXwEwpZtEo
6Pob0jNV10MoQFa5ZznYUTyOz7ZhNxRZiRnDgtahuzvycFt+xNMw7kIWlOFI8SNUbgTB/Hooi0kD
+aCM+SiJi4yxGOaHPI8eNXzV6vZm1ailX07qCpQao8vq0KoYpbEdRWp5cpXDfuYnMHZGjoaa9iMk
jSAC83HuusiWoWs1lAWo+bbrBWXHZEotleBLHEam57cEAheVNad3aXPbAHqYHDtbwfqW/wWqLSA4
jj31+waJd7zyzoIXgjgNBTPvrJEYuQdwaWoWPRip2ejGqArB+RtwgWnTjCloNA0aDtNlFU2xGX2/
tDTpOfs+8cSHiUYHsTLBnR1YS17Ip6OBLXtsU8CF3qbP/Lf56rcmudUYh7mbxwY58JPhmex+Oyve
F938ZyU7LC9kkoGSHlEJfJ82sV3Gr77B1rGQ3Xg97At3tYa1l+OAOdU+DU4+aNF5o83hgMVL/u9f
6WeNCSgMGP5OPRjQuOgteE1j8roIAEFWrUbmSSCUsWVkaGevo+fjhAUi1B0HWL70UpcYqq/hO89m
LtJSGPW9cTE0SDUumahNfgxLDtvui7lD6hI9Ugo5RQPgvaN62TL4CHq7cjuvbqtoL9Z0Wt9frvJN
kgTHggBqfxnP4FosBbosHqrj+4xzkWRNx1pKOT1MHhkT4POd1P9JM6/Qg6MM/R1DXU3MNEGUliX0
/E4hTjkNsVjLvgE6Jcl3Z4W/gC2YKAeMNz5uqCkAI7mhcWExODF0OnD2GkIDGabygohhzsqosPhf
bQmJMKQw8BOMHRCA35EM4OqA0gJC9ef/B1Zo753qVUSo0WeDD1BLX1p/mGGNOXn2FbpsiLsv0tyb
mZTivmAf3S2XhkfRp7UHcuBHQHugHbd5Oi+nPbYHZ1Dt8rFVZtufYBmNEXkgTncHm8vU7Me1ZCup
RsJ/gQfHWG1tOvpVSoRq1xZldvBQe18QSywNsYE26B2YXpcDI9/P4EMJ8y2wrPiv++SAuz7Tc0GJ
qeqLhfJaVpPcm0R/HiSUOHky7kpI36F069WQWpfj/wNbYLZaMQrnbfCMGjQxiQW+bpqCr2IaMLKY
3dZXHUHxygYbuc10s5p2M+VutBsI/N7SgLZJOlXI2YhvtRnyn7sVjQ+isY3Y7AM3R6j6HfzgJW8a
umviHnd2vluoVLdmENLUlxUy4vSSIEFv0iQ6pVqMBtPmWMTpl6JzVh8HIYx2x+OHvYvBQOhSq79O
dBJpfcxp40ZTTOMtu5FmJmGzVxqiX7fS3/gQgBWGpliydQVge+dJ4nXhvnxvJFq1HIdkjEfekZlG
q9v3lMpG7w6+mU2Nne3dRgbCQmMH9PywMPBQy68AVCphSNliuKW+nxbPzk00clf0c3GMfho5yrb4
g75Mb5hMhHV6sZwecfIx9PxgjZGWB1qJKWb4ddj5MUbFjoTzC5Q8oXDcazvitgDAMuqA0k+ASF0v
/2JV6aAhJ6jDZQirC2BcJZrHrigw5v9iAmWWqDUsFCbyRPNy18Y93+XU5o7s8kpeXcdmvhbfCeTn
XDB8rDPM5Mwc2GEP/XgY1JN0MfZKn7Uj1FINQMVSxUKvm2SKcGAShegsVIs5pAW2ngD+GAjzuzTi
PjiWmAxkB88WqeJKU97BnAb95vGk1eiLCvII/zQct+/Lf+iYf3UD/+C3sFPp4FcphKZD329ZzUgz
wcnwWAOghHe7wub5SfHovs5Ia4P4p9htzpgQPgqMNDGywc0EDWEmlekQEkgkHudya7kZuMiP/lxS
Nvws8zdJCLka3gOIeRHYWVPbXm/AFdsN1We6LufJvOdKTsyGbhat/c66wdFU3G6quQA948+uAIXU
vUhh0PQlcbPkgy1J0GF2DLldwZ9lX85r7Ys+ioJQdKLV+NJf/h1u7CmtZboXzXibNPmjlyyURMBw
+TmtbesvvM0IrTw9t0XIaEJ7nXIL20RqSo0omd5z9YhZXQgowOdpwG5skFwr3UPhLIXjc08H+Q3o
iw8hFgPxxQeFjqJDmqMkSaHyVJQiOqgE27suXNmhmVBxBSWi/RXsXESyB3jaqJ+pGgviwoAuM8IS
dPbq3Pgb5UgM1fJkiyKf05o2dxEuH6oI1BXvYlO+qH0uo6Rn8j92P1tW22sWd+COfpLbBIKSos2u
Ll/iqsuhJxWIA7szR2pXHslXRiwnsC+ekm6AzNxxC7hn1OaxJOTDCNFPNV8KsDHfyqr4PEa6zuFA
5ZF8kZxf0Cn1dUkZ1BS8toh2fjhSYLfUZuLoMUXZJWJfOUUfqGJtcJVUyg1PMJbJh8NuOtcX2j5V
kx9aT5wW0UW+ssYX+5G2nDdyfY+Nxx6AnvwVrHh+/HaokGgdsd1dQc41T6vC0KnofWEVppuDvElS
3e3UnUIQ4PVTlAsxNVKDcEpY+XBWO3k0Cj/tkU/5GOwp+dsTDi/VQSS7Dl4KmWj+femRHtmIffkq
13VM06lyTc4bhq4cCpVCJjJ2b25FUC8zRnEv8vbciRhoA0vDXvS+zlrEQynnc4H5CK1ly+CjShX7
d1nfie/eCglwSIYzisBScnqiiQIYt9rxFoY1AhTyKFxf1nnNbdtE+DGkWtnAqliyTTGEtRFFpRGC
yy+8VOCPJn2lRsBr+ZSeuU86+1BTvIO03Spy66KQ1Wq6fK8qYPGwRP94T9wGBbTGRoCdQhjNJ7ul
vAibxg2IWvuhhsPHccVfFlLghuizfvc71zA3AeznJM2OkZdEcEBPZNX4O7cLrak26nhwnIregvVR
n0L74hRuF46MseCmvDh5o8hszO0T+6uIQbTYAjHOqKOrnDKn09s2/d30tH6heXfvidBtqmN3VifJ
ST4Zz0r9OV8JL7tj41mLnIQGXTuyGKIp+M206GhUdTbzrQLrWEzM88QP9R1nC0xoK07D9xIlvkMd
lCuwZ1r343h7a9EPS7X2UC24Z2zjUWA/LaxtjBNGDVWiUxoQwpR1zseMfK3igK8VnNvxdjXfVle3
u7vn5XzNDGqNgJSxugWSf9IyVKzTa/X9c83UUwKBOV1wvYL12iYoJfcr/+vhp/9RW0DKJJNvkHUA
JFYgLCos/8da+4QeZt7xtKTmiSJqoq2YVxXXwEZGFWYnsLFIoUgBVS+LkoBejOd2W0yiD4114PmJ
rjacr+Lj56/hFs4giv3zoetsYL/X7bMC7ZMmahdOgW2NDDtwtwIHupbo69Y3fUmubEpCx5wBdPQv
SNXdVJwObsquqcD7YKkeeeiGSq+05GNzDPMAubDkvBENsKKVkDGMU3JNYyQIHmbWRonWgnttpBH5
HSaPscLPZ2e/AlhXWpw1mvAlBW/B8waOe0c5p9NigDBJvsoEwFJKDhuAuP7yu4Kuk9IzCrIHQOQN
uyc9wvYeZ0dKCkUJJhqjxNgq15dS/bQM6JA+6XtGQvqtac5IQzpKvjOG99bueH/rXaPzlhlEPPqG
6ng/N0PYl/G2Njd9q4UB3/6KIbTyyvRl22nusFyZubgLMvJ7Wi2ijUsL1K7yRrC6fq6ZNrqHBjCR
va+LZGpVz3SovVkHgFDH7Y0QTPPkJZBeg46VwMiThz7RmL+bb9o33zQeQFF3HV0o8+7cFwFTe3u+
4NFdXq5Z0/gr0tHAl+RQOzCTkX5dhFtNU6JrxgDVEwlPxjLetF1W6lUJpdZDTPTY3UogwO5lRmfV
o1pAlu6qU1BMU2yx4j0Y7N6EJ8REnln8M5z/B6Ns6Nlz7eiTQJgxJifgbZcT5vyU5w5HzQB/aS2s
t7uRq57fOO5G4wCHnkz4om9SeCzdKzrtwh/QFvjqsAJlt6M65r3MX10+uJ42AO2SWpyTWOsqztQd
m54l/yz+NT46O4h3anKRF1fdKFDKNym1IXW6ElItaJc1Q2QBCErCQ7sEya4edGzvxuuFi02T41FP
O6ef0iBYp1I3BSEm29AUq49LCTYIk2rIzcni0ua7flYC1Xn0KMmjQxDyU7NVfNfaTyHAb/jglsjO
o6LKnWy3AO9yvbaCEs3IB9PXBY/Oig27ckrFwKuFqKZTSMiynoqo6cvmHP9VoY2toneH2Uckxudc
KDCt4aYoy0zUAV8MMS5WbWhzdMZcUbqFKooYWnBdVLQjGGB/yaEOCcr9FQS92vCl994akl40Mh4r
Qyo600uq9cMgL9aNvH6F7zsCnHDAZvwxIe903IHc6Hf3kkmbPPRq8Q2lR6KdtElUjmY1KYNueqYm
t7s3Lo8bioVS+jZmMwxfu0VLTStZ+5Wp2iTdBhn0C/hmh1B8kiYlzeaKe4dNMHB3dfCoEck2DoAB
LACV13HVbYWYPiuEtKbFt9LukJUngNu6C4PKMT+/sS+hw23ZUk7MM4v39luagLwf2YVcEeJLw/T2
67cxN4AULeVeDZ4wplizQC5+2bwA+GXHxPDPaJYbz3yY/uYzUiWsB3mE8LJKgJ+mK1KmiUfHvMfZ
Rn6x9CKu2lF6suat/sLCx9YopDmvAVOi+gdB4YCI3U27RluOlNG2fpy+fCscX6A8bnFfBo/F1Dgw
NimKu8ix9YcDYGoDDJ3oe60RgGOgK2uVqmcuQDKyqItXEfbYTU/0oUh5WOzr0BxjwD9DI9yX8PfZ
Y9F5HrVgpqUUUmoeP5ZHqRKFGv0GmpklduipujFH1eOPDwPlIF7vRMrztw70C3dT9hbvp0wENNeS
D91j9LyGvGS7CdGsPvVx2h9Zcebgqc8tXSUT1uOSxMVTxP4eNb82Y3rLS6WOscgLTgAgQsJcJlx/
2NHg6S8SSKAgMCUHpqO246VLaYDp6gF4ki0IDP4C+lp80N4jf1BtqKQFs7/hgCbhPvNDr7DQFI7L
f1MQKGn5qdz11/+T6+JytXLXGNsdN6AKppuJ0PGtb+28W/4pO08PSOXg3nM1uSRXBjISPk87oywl
GdrC1KpXZ9rEXaKfdU2BoZCzHprvp9Y24crJvFJ/c+7gTo7m3IJSpEs3NPm/YSMpVpnc+DvKwLgd
LTCShhgAv/TuN+6OE/JyFTV2oO1Wjap2VSaePVYcFf8CXm/ufdYprbv0RLS72YOvTNTvyv+syil8
ijbnH5zP4isS9A9EkufWblF4SFzknlANakgvKDJpzBndMXROhpEjP1UeylcojXSAct9ZyVq7bae6
5xtCy/jaqPnTJ8chNxi6nUTQV3bSEGkCINreZigoWmXIAkutVTrCPV/yVcxEbM42GFJVn0kvJqis
7EqW4kixhfxiPMLXEPch2eiDtG14cYhPuk5gUyuoSh/mmCUCfkAx5i+8TaAzKYZiwsWEGnuRJzDS
zmQoL+WRFZn0UBFfPV3KkWfhimL45Pf8MIWUMJ9TDK0PtiNWrDDnh+1BNU+Oq/X1WyZHSHf6mkkc
iTCotgvH2Ys6lvm75NXYivvD8qeQ3L+d9hdqvApcD2+7sY+V3OTsAkzO72ZIWoO6PE8Pvll+PFEq
Ds3hudfmxwsWd3d/x8x/tQ2EhMzE0LgbWdzk9F9AcEK/r8LotNkyj+NyQuSfkUn64MCSuoUhSXJ4
wJgP/qMWffCUKLUn8v8FymfmZoWNXPW1eaKFYLtsio5dUTlxoYiiFpD/pUIeCyo21sSMWoSHRKC7
3fGfLbj8UwMcwZQoEvddw7zRmhAmCC9RIfxTKBfdURQitS9LXhwF+uFihKgXPtpKfUDfGgrQlKSi
wjg6/SUc92ZJPwaPU7amNrcj1egyQnU1/xFuj5ilLPkae58UTivp5rpjpOfbJjYGkvtA2YXmCshb
w7/414mrEMGB4wEl+GfxJNiQ0Pn4GAY+iN6Um/8GFeP65syjDMHH2iH4eXXFJJz5+XJhc7aH0f11
qmPJRuH/g8fl9iAHxDEQpFo7QsuAr1693QnqkvHuuUhGT3drMDT1fgzza182+16a8gHy8wR+0NF1
/s6I0cYwhdSUluMmDebfRAI75Dn1Dx7LpTFEwzmUqjQf77tvkaQIO6p7UgwjCo4eLW3Yl11VKblt
Vgv/GmWJBon9bRvM0ElTPxt66ZeypLJv1jS1iOIjByMkgTXF/vawxTcKvXQIwejuO6BF79hCDpoV
zQ6jcMRKX0d5S0eGfBTg6jkjYPRsYo8JaA35jCrt3EaovXEdEwpx9Ti1HRgz2g1KUZMllPpXY/I2
op9S/541LtJIf0KhUm75R8xZCzV7GDQKliQQcQI2jfpjvfAwbOM5x2wXbYHMtIqeh9N/9EBSfCQJ
OZRKKobjMsn811A2JIAO8ynylTLoWeHb2TYVQhldPWW6N2pDUEHcpcC7Zve8qIL/Opi+yobu+VXd
TOawIfFzLKCBLoBtrVYTCKQVCBOKM1bqqLZGtPys6uN9n0NvU9gFZ47+Jk3bsZ4fTg0+ujJr80ql
Ee0qeM+TAzFEqUy+YSMMDTTQzDdqC/aKy51v+NkdIDKX+rL5dbbi7/cZRL+HGlpI9W/p4n6iwhyK
Ls/EUl7XYtr8Kd3AMwChQ7rqk14dciAQdgwbxlgXskB3Pi1/IVC/dfxwSXjrKXNxFswjGynymPpO
1lJgbRk8eFqmQd04jQI6m8qfae2yNZmxhq/uOqyQrvEXnIaCC/9DXnKHaxUb4bfU1XbLsVsIs5Gy
pDfBRktAPM95Isx2MReLiIqroVdlj4dKNcbrGZTwTf1ppWtYTFfwsuiNin8AzvrFluW7btAKnZ4t
jVHpf3OouxRV5I2VEKBdIizuzNLY53sZq4lpX9F+BlJzHWUnWvNQtK0W3jYV+pG3i0LypUvo3KYZ
+bU9uZ5hozT37VxeZUksWXThUA45QuomNkW4KnIsPCzt9gYU3Uti6S+QWUso3iYrcebAh4nrpmVn
hOfPDQWQu/T6wLRh32nIWo7spr+9QNn/moGTDM1B0SnhJXasUoAzDRv2aUIhV9+NlhPpf60kwwpv
BemhiHH2LiRAo1V+YF8GN+NxS2LwOZ0nVmO0In8a2qs6iFl6zG9K/8oREzEer+LBONa3dNZVZYZ4
0jbZPNZaRSeER1ASwYHYopmx/AHgNLgktnHbrEq7gji5bhL50HGiWnwju8oKwyq7c3ovYIBCr86f
kfqICd/NYI8FD1NxrI2lTZ7E3vuOIYSZ/Jih9PvKULdHIRf3+f64xuAk7mX9Ud3bl0gsi3ox+U/B
ctN2JN1ww1wSyQNTalEy53l6Bgm/ZvmwcuO41xfuVAfcBfmFMIOJH/Ts9ye2QVXssjRl+dgcVC0L
srpCyBfgVaNCHO8QTBiUxCdoySW2SwEsKhP3cA2s00+FQi048moUEuYuhHlsdKSUkFus/86u2UU1
Q/O4a7J5JI/Mkn2nAjguW7z/O3XgSEAKOkt3TU7JKsHgNR5n0i2Ttz/NfoPgKFDW4iZ2HHpU1I1k
FANUY7iFtoh2A97RqxfsIG0cNARMgNN7/rb9w5BkAb2hflGc+96cMASyHB1zgGyC9zM0tDPP9iZa
MWhwO2fXGKYuByA3dVMuw+2ObAngg79uDPZKcp7dXmLPEKvXBHQkP/plfjfSZBf/aMmy/bmgGtL4
rKtkaG24qJk2IL0xUt2gQn1I3NZIC8csYUufYFK3e0j4Np22/A2pAdgeDH5HNoogTfM74QxCSB68
0Bof+5b2axW6A4vvQgYfzZlBSIdGIk0sewSCMZXYWiDRRM7Jy0rD8UOJqXEpv0tSFhdAlbGoB57z
4RROkCoMKU9dEZ26smR/itWUsOFwF3jIO9U/TVmfxKz7wbi1IPk94LDqlsyhwwssjtl7iQwS254r
eV3PxEh9HgAeAIPB4C6BWMe2Lg2iVLdzJi3BihE6l+q9dPw0Zt4cCO/9slBdBDkkYxGkuH2jFtiq
zepGY24UY+qQJB00Apnthe4Lz/yKhNloFiVE0t/SVaOHejGNbzevtYZ01aOODnFt2P0c0BoYo7kA
IL936p/yLxjeSjUfBl9X7KahlM7JwYBW5JP4NeWaB+/E0h03jtkTUW+nzBWSXc8CtyPi4HWDTDXq
VDC2PzVQTfk/jzXrGTXQP4D6+JL5y7f/iG6i0J4deFj1o2pW3c4dhZnh7ugu3hj8cjQD3EhyYuCu
m3ulZjObqkp3Ff1yOEfPrNFoaFPzVvCFsneag1SfSJp2rcX6Q/myxBLIUDJV1l5MH/ZCGA+fQyUa
JRr7Aa9+B80vu5JCILnhIJ+a2VwdPY9eF7VE6EZSJu0NR2049znOMq1w6ae7YSWMCi0s0IMa0w8e
FepScH+2J3Mc9WycK0qBw6x76mohEisQduZpeNo7B633yLJA32GjzbQfJxxVmQJIIhBgIglhfddu
PB8mgurqILp3mUBBdzJlgIR+FHGHhye4kI6k1ePMnbaz+F83J4yco4cPCB2M7Isio/ljFVU/1lkb
Z92lMGNOmlb7pvUu2BRo74ALLU8PeKVYvxHBykFvssa+5Yt83hK1Cfho93XjeSzKw3L5Bq2zlDx7
re/TQmJslnLPVMqmen975mrSncUOgBkssmP8A6U2I1M+o3plwpMCQ0kY/t1f+msZaFL+igB/fmnL
Aec3d+3jDDjz2ewqaqjkcxtUPAC3WVjyKjYKFfOWdVyY4ei5at1yWiiheyN36HzGtMWzxgUJJv7B
UHI7wlnv2v01KgmcaUF1rFCpJF6cIMftj8MEc95ufZKdtjCv1vS0LdOqeIs3wWUnth1482cw81Vc
hxJ6R79J3IXR3QS6Xi36Fd5WjXn0XBA6b5/BbFzspHCw5ev98n63rWAAH7PVwTLCi0vpLOhdNp7z
zIDakmlLHqdcqZb2G5TyIumZB1mLjR/z20oDezH3wTmzx2y+/nEJAbFXs08jPanSchMM8hsBXO9e
yhhY2ndIGiQkzO3vjylBAlCPdy+OOejPqKnTxxyitF8lHb3NX7SnyiUbg9cJ9a+rT3AGNv7hf8z6
Zw8vHl74Gz5dJTCXOmtYydSHAX3UbNr39Jh3LTCWbyo/nDRcwj9hrmGw6kwuVv0ORP/AxOw+yk+u
HW5GAX96ZEfF5XySgjCC1wUeJqUU/S2t6NIND9EsZmUY1X1+6PaAsiAulMmDE/ofWswDgar2fNiv
EQhUjKpp8AcK84qbLl9rIEc3QwNTW7Fvjax73TR5QOXpF+27dzXvlkjpgOG9u8zDM5h+psWaTAa5
xz3rWY5eVXRDF0pAEpEDCCZ95hwT04BWi5NgeUAGUUTPqlBDcc9vfnuTvXMeBVwPRzHXehl4W4O/
po0vQabW5g7DTrVPixOj3MzJOIDA1O9XFOHn491xB2wNcArUbk4x1faMSAcRszI3x79D1q7gjuBb
WHzKH9oEKW4OwF2ls5EthRMTT9Vl+fE9WAFLmLpV9WUZV/vip+0hXriZBjp0kCxmQvJheIHtN5Zy
OYqZXm9jp34hDbO+wG/TLCNf90hI05rO86A5fkpEytC/wr6vUYSG7t6zuOSlifhUsRFo6XqioZ14
nWylj7EMNuKUT/EAc/tZbqJWKOXEw2SFc+wMe7F7h76paFhbjQa/u3g2aIcSCwKwSoeTGpOido7a
TrGA1v1oOjP2QsZKcU+d150WHefTb63I+W4UNSYqNNmCV5oCGYY4G6tQlXrU4es3omCUHTI94U5f
glghjz9mWWLomFVobrH1HrORTSZmQ10TdX1o//xMNVMAxVBRd6fcfwYXUGxqyrspBBxnhPztcALo
iu1lbD2PAM7y9mFBic8SA+NfNdyxgb0cQ0ixP7YqzI62fM3/RB1r5YSfI1NAg8eTbciCBgO2FtR0
++PXNrAFKa/5ZbbRGvqJ/dutkiHk1wKKjm6D7fkZuNoJmeDGH9Iz5nrz3Qd7E6lgEuMD4ZnY47lg
yBAiOSRPlypZZI8ozrb/h6+peTOmTk6WwWDLFrrHOLMY/nqP9blXac2f4Yr+Dtbq5tGsh5cRp7Vp
l8puaEqr+oec13k6bhhJIqvBzYPkVdR10sCG1EdJQmkZpCG2RNFM1fSAIr361DAlWsa8LYlJiiFF
JSGnYq0FE0CeAqnbynnNHWILFr8+W/rIEGvXa57c7deOArlpXBHtvFNf2SGG7ixA9Gq3hN3R2Ed7
l6M1CzbupL6kt0IVR5i8AOL0dk8KiPOI9+U++ijS89WfiTu7y440ZJ2f7nPjjG0tg3tKepDp8MM6
qD+/ng6GSbEV2oHxnDdSV79r8tzeX21V8ZAq5QSXXpHBOPvaIv2j0+pnI8s883TV+s2Fcv1Neg2t
DzKQ43x18/NQ6VVzH4v+EzAdKpEpuimI+cHpPV3RBmff9uyrwhwcWdMgOiJZF8NQJVKKEXNMR8OF
EVP7HlrzvKiOfipdz8GuSFHV7tZZNrL6Hl99/WXkfgcutw3f9MI93wpUrgj1kOEuestiRnf1cswh
s5/9eagACzUHFD02LqiclFlBtWH+gA+tLxKdme5TKH2mU0srmXwuAwhWqbqPqykYRqcg006hhQIH
bEYs02cNuPFlazEBpCAtnxm3Q98l4iVD/8P0lqVZIxKencjFTZcYCgbaIl4KQS0IIexAi9REzhj4
iCrYS9d++SS4n56rHH0tyMaXHX2q7SYDbxgE/XjwgNBRYatpinF8aO+o1Z9qkcEpOlGpCi4DoWIA
xeFe3URJKTDbukDQeGqyf1HuHAdsk4I2rTG70weH1g2ddZ4POfhhsoI5ZAtjPGWID79RzH2VfZn8
hRvOfXZw6LcbGzGUD1MFe50Jwvcqi+YquMy/+NH1jXPy2aZeYCseo1VnIL+6pbalhdl7sBTJLa0J
GDaEgvcHcvnGdQeRsjEqELe9GGZEIaTZzS6Z81O1t+R4Eqf1akntBlWieKTnDfX73eOhV3GiBp5q
cvuHzvGhBN8qGAyglvMNHzZjGZ7Sx2RPL9VxtcCtPMW3wkxETlxQsIV9MKvggojb3eh2uFRPTKpa
fAS0qwvjUe3YN3OrwhUOSlVeeZKurm2qRCNEnFvxINudea1hvP3Sqx8L8fWHVlxaRfLUSb3BBZIP
5NdktfQ8LGGE0Egq1g2kDrjbozp9Ms27vBLQco7n+TEuUAixOIbBdfnooEqUU5wPtroB6RykJnmn
HQc5UGVdLww5tWO0gxCNTmHoSPQx27Wb2V5DmYkT5em8ExO8UCSSWhTnlxqXwnq8R5g6gsuxPrYd
ZR2WDVP45qooJ7LIg7m0WCT1FdQpdnk/r/3qbmTVGphd+i+KRDvmyIVDz1DpAXe2FXKAwFL7aFK/
ZVRf6oDFu7vCWqikk6mZ8zJSfVtDRdH0fD5SJrIkDGilRKYesviZ4c3oKYhRNXTqCIn2Hewcbzdp
KVBNcR24lV/6lt2mgQe/lzfo8u1wTYu7bre9IVtYT4CFBa3sPAG8eU4j9uQubnaFRH0hynzgsiCh
9Jb/yMfR0PkT+uMrg5l270mJxZhsqBpQC6qZNcfgTC2haSq3YfBYjrEhy/31pOOjCa6PSQHHkW9a
N4ccdnwdanDWZBraaLoosCeI7+vKCeEw6DYB/8bqoDh2ThhZXVV2J8NZruTKZ4BLVmHJ9Tgx6r76
k2qCDjSM7y5AjBp+NJ+llR4PBy5cFKLT3a8NNHRVAohShIHIaemxE7ApKNWFts1H25DO5BSGcQGE
TscDDJWSnO6tXDtD/UKu61i2MTycml/dosp15gkIFUIfmK1ZfpK5OiPPLO4amr+p/czIjuOUSS8Y
oUZHtPaDZuQUhV0iViXsVrgJAkcDq974PIwg81Zod/kU+FbGgGiBQx/vddnd7JF4mqINNURPL+kF
k285dqDUwH2viPtptCd7BiqouCpp8CJJxz6EXbd966l+yMLydvcmDs0qJ7t6mkpRsFYz0QMDDnnR
pmwQV/AxsFFt+oOr1AYgW2JWCwJP9Az42SPtWDVWkXNGw4LkXM2FQ6BkLZDje3seCSF3Ns+BAkFI
JmjgtT4r/wOtwdrZG6Z5pW6t0F9p10W6TKdwg/emajJtx+hKKpU7PjPDGEaOnOlcv4KVMRQt8Koe
uUfIOD2mc9Y65ZtffItOsoRd3Goiqr7pHhW37IYxt9W7+GXZ7JyumPlw4D3gnwiTnN19s6O42u6e
1Yxb1rbb0zDGO2scoDvQnmDYLNhHyzWbYjHUsNd2sXcVC9pJREQMsCzYuXGuYlhxw9p19zQbU1So
s51leT9Rh/fH58ZkkiLww5qtDSbFw++cT39Oq96AuilUsOlaQLk9LcCZ2xmNgDeilmntWnOZAolC
xfiW50U7eO3FIulFAgwzYN0qQTQ3+T/RGySQ7ejazgc2wU1qUAwWNMgnkKbwWjqZW73/QJ5AEFaZ
/bjMkx8so4uNCWepEcgvgVNfPjKJeklWIGlTyz8KJqQtMHmedHWF+kGPgMVMa1NkjZeChbKxBJMu
t6I+umzTMRxkT39ERbGWvGOcAkfezdjha3xBJjkvTo3orsTPVpTaGWPWPFCdd9I8OaLLuzoLjIXc
zNOSRs2eL0A5rWAXunVEt76X9JYsn/2rOqO5/CEEa06oNSwALQ9H3/6i+Zc7AMgtOvyTz161AIBz
qIF0wRGw2kmNe65hX4uqQQ/29UFchsQgrB6M/z+3b3p3eWVLjQCiZKYnFi6BVXJZWnF1PNiO4z4P
SBMCsA7RAV1H07fpFuHiAv9lqGUToI6JAod/TSattlcS/FwVZ3DVLxY4HjpwDD5RYvrkh7rTfzXN
CFAxWfyCntQK3b+1BgKht2Z4luu8eupFFd3amp2FZpe8L6ZoR20QAJqfhntuCrTO2zk15pis9HLT
C1j/3WFg4NEk1xdZJsOqFCR/Te9tuZeIjojUIODfxtTt5LCAD1ATrC0Uv1TF209MNh8RBfWrGkV+
hTkKPeID4GZMddJXpNYlLis4uI0494di9kOKAug6lYLBhyOQA0Yhvs1pEbi5Ic/FgwC/SJ2r0Ffz
xHDiwUVcPCBVQ6wjfUHRwmUVpPa11RDNaHGuoQrtu6gwwS3zCOmxM0dpSTUiVq0LyyFDeyTBpqRK
2yZZ3e/NV0CtDAlKaLQ8qVeqQokmaJRgVZZulPF3FUBImunCn3wVPLpzVRRtefktFXX2pcquuB2/
jaODHwQaxuPeZrReoPEOrERwNezNnAfO/GQ6oynaxjWAu+fv3++rr82j/G+kLu6cl5HywPHmdcNX
UtESoPzZqURxAsf5H07Oo6ju//86jAbBZJYTlQMCQbrcBQEy63rZqoph1Qfydb3he91tCSPcRmCb
WeaZu0zoplNUXnoDzcbMoIpkB//axjaI9+wd+5+/ZYLsjczJxhQFbytMa6ii6ZkIceJDkMv+HVr4
CynLXq0TruN78z3TXWt5DHsbSIZzMWfN4A/FsceX6JWvgEce2ijzm1AEhV1xEfNdnmf4G8x9sz5i
aiC3Cl2vgw5hY1cIj1YXF0HMhxWCSVd2ZD/GM+NFwsTxplWwP7t8DObry7cH5cDEMXEe1wFxhwxz
sDSopGW2vfLbtDH7dSuLddnA7U59PjhRqOzYsas2YpU0LsRgQ982N2NOqp44H97ezn97LZ5AHUfl
HO0QaV8l938qYQOLd4iTtrD/LLNWV0ooV/Qg0on9eMVPf0IPug6DvizqMhathYSy64KsGsh4eJXj
lDAoN4MH/y6ObdjKgVlEMpFw+xWPzA/MB097kcXQB6FnlRCYedv1yyP+vX/G8VUKWks5XabBEMlu
OomjYKQggZg3t436xdaIUyGHW9kewdKSde72LhqjNXa62Yiz/XHQ1CYCwpgsOpBuMDL8K1oGNpEJ
qIxGvkyHzcMPL6ulrdwmn6MUM1P+0LpnMw1MR/C7pVa+LwUTK0IO7gnCpr4zMfr20v7kdwQjEUNK
1TLCryo19wJnwZjJRbhCL5Jbyz3dCSWx9JE6J5ZQQNu1Ggx86PsAUV2pUhm/1iJAVhFirQvN8yDh
i6XumS+V/UsnZOxnYeBN7P0mTuP7Ah7yaRBmkpGoBbgwduph+ZjeVuB+hTGEZ/siCdNRXxahjJUD
z6af7sAgDb+addnVgNeI+R55BVgxmym3Pv2pdcdUH8ZJ3RpXNalb/DsTwa8joFWp1ssepmOPvZJZ
KWRwRGmEyJ4Ac1r68t7UhWdlI3+XKh6FuKColKUEDLecUlZLAAlLwLYQwliwLYJeOLVt/FVej63c
pTRTVJANZH5vkqvfiU/5cbFtCL6yvh81ZpfggovYq/72PLM4CFbUqJRfMOFIC743U8YgqfOLv4lG
YT4pqZTrzKeV9nl44wmGUwKs5SGZru3zBhwWPeOwqJOkoflPwyCaw+i5mX/Pd3nTdBtXCl3YgE5M
Asihampa8jpSTIVRXUce6rI0VvWz6l4dCX6aVvotB1eZtjTg5ul5GYTDYdISpfwQnJyIOazc0VrA
Nr1LMPEhWelfKC9Ha1spkwk+2VyO70LUQAxSXm5oVDeSu2U6yEwP+nnnpYHFaCKfHFEj3FX30O2O
hp1Fj4v50y6+ot4Ivf+gOk83AMiWubJjVFkFQpyFYbn+qkH7ZnjEPlXg+8aeTY+Tjbt/mj2EBY4a
l3mF5H3lI5FldDbQkifxkaVafQM2nex7aGbsxRuRcrfTB/JxZbWdTifL5YTppervzw8Pkq4qgdvA
YT3yUPpqw0mzp/Zmr/rlTI0MuoRvW3LkruunWAuaD/YTDsaLm80BdzG7i1fY7n+IWr/BAEBCPzU6
tsr0+KXtIe9Q3Z+mkU7rVKkfd66HkdHGKQeqNCdMMLnGeE8MJYqq5tUuS4e6IOm49wniZNct7ERL
z2brCyhi3B1Kri+eqN/sFTGDIWI1fU00zPtlIv4HrS4Gg0x9Uu8qxsqSUavbQ2uUC8e05t6jY2lh
+f4Eun39Zz4Er8yRD5uyh+4opsXe2ArMKLyLVBKeDeMuZXML+CKqa4lAw4gAEX0NlB+daxpAZKtj
J0cVaBPqNWXrxOsB1ZqpxbdF9Y/ydI55jlJnDv5G90wJKjGKElt+fKb5o65b7TVXBzBPvcNiLEct
bDGZMgZZ/HT9wGeJobmUjsXUoLu8+CVuBz97B9HuGR1tRMgnNUbOINTnZiQjy5BZZFSMMhbI5HBb
7WvBDA2WBUNIuStSTHe40vIZTXwUVVJO43Ugq2UtOGLx4gfC2JSvB4nUuzlQVPavbHnYf7pz9CVz
MPK/7i5SyC84AHgUdQtGiRh8JVYa2ltBV8c6JjG9hfq8jqlik4OtnQ/NdNKjsjcxBaZ3OmlWfjfA
IoHE1XkhIfJKBXRDFo4x1bBRXbTq5I13ucl9nJkGNBpEZRdb/5pRFnTx0ESiEsYlpKbmj7KAoT3b
SBNyHN2jlbz7faDGC8ZxSE2mRYrBdHiC+/YDIqqFWvaNEoKr21FHDt5mfjeRnstGTDq3YXJpFpDD
qxVw9g+dAx8IMSfl7avgokjOO+EgeN4lWREGFkSMxhoV29WsTIccZXKctX2G8vTLS8NEtP9sRNOa
C6CqrAHT1no7MrgJ++Pd/DHGXndp7EjplZaV+okkd4izZA4+OIj3GN4z4S0VLtjV4VysTjMAHL6P
GScKTT4Xw8RC5NWUqj/2CPhKSqptTL4Cv4i/wrRbN9aMWaPDX9mslRzF/d4izL4taJ2kDMqYtoly
Qvxt5XYIiwauvMfJP1s9R5n5fIHnYF3kPi4tQranj4skplu7QfbeBYbK4f8Zxxd8+wxj/qJEMmfI
V+Xuq77iBYe8tnHXm/4gSiay8lyAplXf5n7UPJ5cyLf7fRZx2l0E9AIlhKX6wygBS9fhMthXhU7J
dbCezhzgUfWMIofqTdg+O3BgqrSe3N5T3lsBP7xQWIMVyLAPoHz8tFZv7UIWeqWCEjzqYDhZz+GZ
aUYW13y3+sYLL1HiDzQY7hvUe9UIjjGFyV7wW7/zZyLo5H/V/k2PQd1xJQq3etdqNu++8ec8QlTj
Nhqm8djf+cU3TXHSVx0Iep74WRWuqoSlR8xrt414/yfUpI+KKVE5jITOU4vMKvVrzrfSdsUWePsE
rnt7kSKoy/EcerwcylbnSRnRZmfZEKLayhrkQc2pOTZJAMDI4gn1oPDUQYvAqZuLbeBKyY8JRmST
gd9enoRI4qHYcHOYAKWUfYuAM+7muP2sxOHgeesm52DVwyiJCMiGi0pDZBBfnEEPpb6UU4CEkYn0
9Q4akI5WSvhzoLvT8n5IAmv86226XUM6oWTFdyuYXbc089e+uI2wq1XGLDlN6tgL3oyK8EKgRe09
C6mQPZr9DQnwpfc8xl0OJneaNjhBEtDo1L0b5b79l2aTVN68BrWb1cCxZaJxSwzl3w6QBNLqFLNW
XjvJR16ac993KcrGFAYUXHAfUfNyi108VO7xojByvflkdsLAolLOzoEJK1/AEpe8hjW/GHrxNH8y
Tj1aHrRAhGg+bgkpjJagvU8qDaDSwD/N1CT8FU34yAWsY4oT1cv9ymIV2iHgfv56rcJlwjkQxv5L
cFfaI/U77zjHB1GxPAiNEc0TW0TWc2auYpPkMJEZPJXN9OTh3bh5iI9bCWmhNagcLvay4rcuJs9f
+Vvs9VV7rsghyxysN6HfNrReaRyKa0dWwDIfXcc31IAaD6TAXv10ABIXVK/Y5gy9LEcCo821PyX3
+UUlTX7PmXWlHH3bLltzdIJ+ooSOGFyJrPyPdDgJbaO0jEU0WsJhOe2BFvUfV26sEFPKs9qJk5Ip
5RGm+YrDeWQzLAkVj1Di34VVramm2RySxhv1JMjVsnTt7Zts7D8Rnuy1c+UM8x9fSGDfHsLYDoxm
GR4LHmFodKU8bC/Ezz9NZfQSmYT82x7OwfMS4gHERDDDgZF346mCMgD3hULNkUwuR6fnlpvVpFty
tDr8670gJ6tAqTqnVoa/95SF3FgAFrxrorKRb8ANYKUpBaEMLQg+Wmf29R7V1eBX+NKdAB9C9TnG
2Z5tmGLctFVsmFzFWj696mYNb5tpTONpMvavCj0ws7W/QFJOmBl1/9/B08yuukZpi4WtTSdjgUuO
Jui04yJbc1BvfQIw7xXkAln1ATpuTSoM9GFj4D4Pr0o2NkwEgTckukXVV0J9BpNdy48lKWPlSm/E
XZey8711zbKL8AoiLlAKp86RJ1f8sjZxugvWzaK2dunV5iSwfhYrddFf1JG1uqwb/ticQ0gejx4J
OSrsCDOSAoGZHz269Q03AhyTwr/FA3pNVnmuIbKkdgMrAfUFoZGZ6hTOwfFMYXQ+UiFLlitoa9za
4VO49E2u4Cukarkp8orJCIhKfu7yyjZotudr85p/k2qebszRbwOiEJZkfDy2So+v4xj/9aPdfCzk
bnYJkYYwl/JRsvTlbKwjoVcqV4z+za0qr7hdKU/98IXTO5MhuN/RWOjoba873W69qxI4SiOiks/P
d9Urh06aE7uZW2zFMl19QPfKa/nshu18jeAP8TOKegWGNMk69N8FviAl8GzWlfs+1gm1ZTYU2LaG
HFxpFuyZzK4/ApXcwWJNKbQHpfk8jXMSBqLAmCMRzC5f/znmy2QI4vXt8NdS/5rVAMsCnTwYyzt3
0N28XZAuMSCGKcaqt/EINqJwG1Twsa5lcg6JiruzkBHhkBMkuc8J7f7JIXLn/XYdyUcu5+pl0WRr
DIGrS664qZ8OEwEhUrBjrD/xntQy1Plw2Bu1NDBWwgicsfW6GB8YuSOn3dzwQbHcpst5DT9aPpnF
GHE7z628SJ+3cmZfuiUgle3vZtlQIiTGmprad/dDQZNbJXe5cYJdhN8pwHOwhLBmDquVaz+6vSBv
f5Sa6HNusT4n6AvnSkgaRJZOBjBEHtnKflOj7H1DxM4vXuvT07eJcEamf0GTDs4D2qKrRYFIa8s4
rIFSfFkbhO2zr9mZtRcGlx+ZTocrOsPdwteSnDdog1M0xEGTA/4w9lrKXGgI1M170M4YAbA+uk16
ju+JOZr+Hh3bqlgJEefYkj6Vr9eDQl2raEjwH4cCLuWhNfHHAt3X59wMSakRdilGjukb72mWf8cm
lZ5Q4GrQflBWpBDTNTBQuGlw+r+GyYIZTmxZVfv7eNg9wCa2yfkZgNHii0aoH7WWzDc9XwGrKz+Z
lyNvwIqaGO5bqUNmOsfdcyNrHN6Pghqp5/dgayqjuI7IospVC8GpNryAXDxLQqhl1hhaeHeqy3YN
Ke4x7n78mtfnGJy/SyuhgVY+AtzxrEvAlutXpvmvZXCANQOcpHNIphmLpCuEvOuqZm8dYowjfc2u
P2wVhGZCvSoVI59pTbsMR8DPyRgRyZT45KT33we+9Q7/cFSooZeL/ECUdajeGTZu7jrt3IPukgCW
qdAHFrtFtiPWSjgB4CGzlrPv58h0lMWWA7ZgkihX15V0kLBy2bMgq5gTcCiwlQcOeTf+1YZQEL7V
kZtj2UXEQqjcsTjVFltXpEAtdpCo83c+CCGskw2hRWJrIL84GXbXTlgtyM/pHjgzmbTPBMPn/X0h
kDDZv5QB4Wlrs3TyER13XA1aU7IH7glm7lRQK9b4tWgMR4fevSTnl9Q1vLoOi/z4KJLd9SDHf4/8
14euOoVWZXnaeaIRuDG9uz7YkSeDRMc+/mToAm/7Dtnbn3KgYlwnDJ9f8TlLAYoLoMXLDCmiexTh
A9pR8mUAM6jO+MuDoOKYfNkb6FjLQZLEYk+F3wBgXuBTe1++d6/Wdyw24VFBY4aDFz2t+VgNlSiG
r/H7AAz8bPF7/08fmlBzrLT8yTUzUKycCO5XsDTwyTemHVqEs3pV3uNZ63norY0bdaK6Y0pwHD2U
1uL7YMtH/l+SIoVt+lnRpiH3L9V9PSP1HwvPpmRFyibjeifGPkxFlB3zC4LPMO5XEVTydWFEXRr8
dekBN4G02v/PZtl528t+MWXqUUSNCvoYw/ZzqjwEQYGvk1Ov0sKZb1vLb/z09RDDMBm/pgRynxVK
pRTScL90rhSrEd/qYQO6ng13JaKejsuBcAhUVfWTygT/LUe9hHbA/+NLoxzndcxi9zg4P4OHy3tX
Q4Rpz4zE5ZdolOD/S5DLWX3qVfLfCq9X30vN6uI/qzjGWbHZnQteYckfs9C9L1jo/v+hr13CbxnM
8y/vnEKTAnMWrchpj3Vo/WjnELWqevw73J2k2cOTD1/oNq/Qq//NquctPINdBfLzh1QxiiYRz84r
yVpxPiB2lLHef6QPViy+O2x6jSrPxf4zsDJwtjCYXPzvbXC2cNmoSNbOJfVn3PVcQzowliv0Oq/F
v+6Mz6vlQPPnGCvyQR6/Du7yjueV6zQgUj4jdjPmKrtmOsBpeCosFOQ9h/81KzG1dTeujRARX0kU
frqgA3Td317XjnQm2N8i32CA9j35NGAugpH4O3DUFPvtCqlklr21IhbuMFj6enoi+c7AGGit8G9+
cIRP2bc+xrfu6FUOfhmeyUVUL0kRfw5omzwj0BGVwYBpz9IS1s+VfpOogp0Ep2Lk2dB7aXxcNMQs
AJDtQrOG9pouenhRUkZHrCZv60SJdxMh2gjTPbRaIMJt67iVgagD262euSyzr5EjxD2GJC+2lCLK
mAc5rksdiXSAERsbhDC8VsMFlJclROukHCzGc6LPMrBVtKOD/beP4Q/+Ud1JqlhQjHt8kZ71zg9O
NCaCRcY0SI7000BND0arkjSeGzCPzPwjWFy/KkBu4gpmio/8hPjtMfYbDAKfX1/TeyVXFSSTDONS
HXYspnInSYq2n5trCd4zky4tAxBaixsSHm5uCQv7fy7rFxn2P843KlOaBfAaMJEkMvqDJK3G3Tfd
I/sqDGnId+Temw8kynY96UPcm0RGkEzgO0NTTd4iHFHWlURpVg2XAnGzEkjUbfxqIcAyZtq14Wc7
jbxdeQpgVmDe6r1TqzzM8jqJ9IL1SpfKA46E7hRcSujU6R1YlDpmHeDfXeCXjGaaMNpnBbw4CjtB
0jfdsmLW3hvgdxU7+gg4IRW3A0uWqRMma/mx8WIoKq4lCPSFn5hBbOTqc0LsE2EBiEbh7LkgdeWA
CdnqaxlR4KUA+jdmlR4xywsRfX0yFKJUCnqaibhC0QMPxZklyCosBDMlgMPvLH0F+0YaLN7SJqT4
A81RpyHXK6B1U+WPh0iPIw+gNcYfI0WK1niECyuqnIcu5WBApPq7HKg67yp9/M7Rsm0aZN9KenYy
ne3GEPmzoduGXr2/8IdpEFtBaTBF16Xqs29Xn1k7egeqVGq7J6zc20WVAgKka9E0zu67lV+ARsPE
xvb67MsFSquce2Y3fZm97IFMsm3J6wqIEI35KzpImfOzqw9X7Ii6oT+uUES2NDI14h+puvIaeL6k
wn+jtn2XgTo1Fpp+xYdkmo6a0orFLoHXgYaz02a1xHzqfevHWx527miS6NInDOzFyeXn3r/X7+fK
nU2SaA2Kpn2zwW74bK1dPmdyQS3tCq5wk06qsHwQiJL3WJCZVAU2eKtk6WCqX7K1QqBrNmh32KsI
hIvgWsdPO8ajOFuOnhdr2nuCEBao9H3mRSP6qWbHzvw2vXOxw48tEe3baAhEqPg9stNkCiqYK3VS
8siIy61TYcTHLtPBp6Sy7V1nil0AP0vkW7R5OhMqgSLhY9AP7Z9phvyqrnk8rp+FmNKMLLBVIrdM
51h00Xukt2FJkKslNPs4+t5SiA0rigtssvze9Ty2ig8BV8zLIAmcZ79CBk1++drN/B3TYwxML+fh
pqAoxISmpxTs9liQsWSHQ94MCKv0zFKxsfKP/NhCUlJrZvsh/rNyXGTq+aCswJl3Q+3VscGrMNmG
79yNwHGGlyRriXpIhkIjmtYgcSfObwBkWNRDxDU95j7aqp7UN3159PAVwSiVWc3yHvLQsvBkkYq4
Hpe2IFfQmM27tPJo2rOLucLQM6q4bEnB3oIxF6oPI2yxD030wc+4vsyMoH8h/Mw008emrKwCiKTf
aTCk56qzIFhV8zBCtK5SFyIhu9+9RCRzNYybzcxmKD+5Z53KQ217EtXvgRa83PoWeIkiobyJ4o8c
wL/fz7k+hSIVlb0YrSi+C6DI4hIqb/YLsao/IY1eeHK8ztYqH7jLnJBOtLNyQOOquZfR3EK7TRBO
0T5e7T+SgMNvdrP/Yoq5VK5DYaHkhOhCx/YL7rtYebF9FD4ttLVEwdHjW9iF5wQv8OjiKzX/qK+B
6Z1Fpg2d3iZgQXCzDDYqGn0NtEc+HLBjtZ30nARSSbO334evr+iZh/lshIHp77a/gqLkqZa0Po6S
PM9HFajEAne1xZ1DKyAJpCgFL1t6+EPLrw1yR+uQWS2tFU29cgapo8RL/WJqKqn0xe/bdEqPWta8
4WMgRfwFlSILP3xl/1ffjrJVQTgzyTb7skDxEzCkDIlYpp+MoKr91lgdgMDqfn9ex3ulpy7Tetpt
T8rzBosu4a3tUXfAAtb+NF5Mx42rqNaPMmF0iAMqOz8i55Zeqw7woLfV4INKUp5IIB7ztv5zGBPJ
NQ3awWdkJEx2WlnCBl/23/tBtEECnTgHmwGedeoPpqRUrK+2Ww6bV6VGVr1V1CAky4eIb/lJCCYr
RHw6RMRt+i1xSSLDVT0/onrBYO9nUNcyEU7oSY+WftzdDUdFvdqzjSI9LW+7TsyZqCXKPeFu9aba
hRmke03LkHmTUKqNyn8Or3YefblTR9rCAy/w/nDrhG3EwgrAb8/I0G26YT7gVy7hxCp3jCoOQ+0S
xr06aXHOjE29qwC518AMBZK69rkLiYOz+cBFD6zapkimJBTiLnRQppRXC9s9phBG4ldF61iAHq6o
hAcPhS8uGIe6eaKJoc1dfyyR3PGzNRaAzvr78IMki4AY4S0oHexzHNdzUeCMDcjcrdbFzmMKZTYJ
lCI+Ojn45auFh4P9IalsRJ1lQ/2ywZSDkBMtvh5vhjHbqMFVcr976CRFzZdODvOhpgu5denKgyDL
KwvZaWbAgbjP5XNlkNfh7o2B1jO8EeDpFYBDf+/6ApmfMrlE0obyKlnauMOXoBj58f1rqss9hkRg
GdBybsyOMukh0IPpMym+7fqkMqa2BTe6L8Szs61DlRmUrb5DVxgUhVZS81QmLpIAkN9Kyfe0sMxj
KeuUIvni8Q7C5Wqj5EkYcy2EUzDHiEcOS+A6OqqNuFUz43bBbgIPfF4qkDVoVMV6h/EnB5HW1RLz
FUCP//AftyBw86wbaL2220XQQTTtOfPSnkxHItt6wbl8QXF+xb/xhM+NNG2F0jFmD2aoSvQZYnUj
3HHDRyWuoLmoI9u3pN4QuxcO4OlDOKVgmYbwcRvBGG75xexaMbHvyvjvEGdWDpWUYvumgSE2+xs6
4FOYrHMlDIu2feANXj/Z+T09zN3w1/N85YodwEpetivq0vYTliond2WbStav7wmAborjBAqhMgaF
CA4ILTxAfqilu883VWxZaIeCDbyNlX+MKSpKs6dplt5CD9Ll5iE5yDkcN71lNKgjRyfdUZhx15g2
Ph1CIpINOEZLl1wIrqbN80VghusYSLWmLsPgkK1hpmuTns67KmOoepICvicBXi8rPV1TQsumD3E1
KeKJs7JKOg3Q1LiJiXdIrwVXikmddGsz9FhID/a1uvyAGNX0iYkh3H9I0caaAZRGQXmFz5o3EW07
TPFcoLU5QP80hSflzK2qYq1c6pTKy36huSlzyfhwdEY02efmOChknjX+Ec03BdON7pzmTcSYJGQb
x93k14m4VLFJynhR1Bi2SGXSm3GI8ZAfbuDCRNdmLVOqk392yu/p5WHOjtma/sG2ybNkF4ln/ouC
UjQT2xsgUjxZOfvBYWyNmvnJnXY1i2DyusSnQ1oLHmnuKQpy/ou4NvpjLB0RGcbhOtvFRzVuLW5S
64aMfchOykY1IBzCefgfQNJpCIKeCIKzr3EXHxLJf4Og7sMxUvHSZrrebfboA9GSgm2nnypQYm5A
ibO+uW/DaFL7oF7iEvay1sgk3IiWU2FMBvXnQdYF0126fOkOd8M8lSvJ+5BztYH5e0zY25tEQz9T
lmRK2gqTMRw4c2nMf6P3BDv89raLVAM17st2ChkxM2GSx6jdmHfAYPOKRcrpL/PXF4Phe9F3n69c
eqkEpp2OSRKwtuAv/fWVABNCVIrrJ4A84vgxU1NZb2jDrBFtkwi0LmANy2UtySgQo+dCkS9as96n
XOVPahj4yz5A+duGJm/8y5GeSNtgFDPvyYHGFhxhl0ZPMbOlH24cqof8kD7+PMLL+ombIhbl5sRD
3ozfKBUTMHt1BcLrojWubnEGlNvpohmWxbR5DRktAyBM0KREi16ybxClwH7JYco4/mE+n+Fd9pRx
VuoLESEcdy7uV7Un1joUYaI2+v5gpiwqg2BlFj7x4F2xplbqt/qqRMzNORtWIurPG0uEA2OYsfv7
OiDbd9QSGNO3iNhuUpn1u5+KT9hMONXkv51K58cdaMvmmtAZnWZjXadOFVhS/6/kMT7i4yUZua1t
q9kvHQmZwzIz6e4JoCcHyWKUw9mADGVwFC4L7mSZA6dgQaGZkIPdtwt6aoOuWTICc9jMAUs1DmGA
r3blHtOR3H8dt91hv6emAdRwYIcSUpYAHujfmKgl4dlc8nGH2Qnt+dpa9EtCamGzNOLXAPdCi6Dj
45AHf0b2YVjw0D3/8+CuQE3Tnauj3nz+QYAFJ1NFf83P3CkKZqIW3lqdThqEutpXA6IDxSo64i6J
CdLx3CS0MF+v32tora+2B+6xrTOjDSwpxbssH402PPer2De8GBKHUtKCFxvEia9i5mAeayf9fq7H
LN6WP/397UcX+cGfpOAwAJiHgKvwM/7KNiRs3cQNlNpvf5s//cgaCYUCZQxiD+BjdI9so+Bj47UI
R832SxCr420qzkQZI/gCl0IDVILbnE/V8zqRJZoiYQCyP1aMtmCP7qmvpaUYbs0ocP36Rb5K3LLS
aAPSQS59FGO0nphWdXzO6G1/7hJ8mc3n2FNm3hIKgXEGebqHBfiKyGDQV9PGWoZ5Hg7LdQhWviuu
WhmZIl1vyz4iQ2U4YcS4n16uuTb3u3OlJyEFmFYFQLvv8azn2+MwVtAdXVKXHHTn6/PN7cDCdxb2
xK8IWQ8igh5yVvpVYRkU/suIHbzdygxle7tA2j5SVocxiervTe3p
`protect end_protected
